library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
ENTITY j6_prom IS
PORT
(
	address         : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
	clock           : IN STD_LOGIC  := '1';
	q               : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
);
END j6_prom; 
ARCHITECTURE SYN OF j6_prom IS	
signal qq : STD_LOGIC_VECTOR (3 DOWNTO 0);
begin
q<=qq;
PROCESS (address)
begin
CASE address IS 
	when "000000000" => qq <= "1000"; -- 0x000
	when "000000001" => qq <= "0000"; -- 0x001
	when "000000010" => qq <= "1100"; -- 0x002
	when "000000011" => qq <= "0000"; -- 0x003
	when "000000100" => qq <= "1101"; -- 0x004
	when "000000101" => qq <= "0111"; -- 0x005
	when "000000110" => qq <= "1101"; -- 0x006
	when "000000111" => qq <= "0111"; -- 0x007
	when "000001000" => qq <= "1100"; -- 0x008
	when "000001001" => qq <= "0000"; -- 0x009
	when "000001010" => qq <= "1101"; -- 0x00a
	when "000001011" => qq <= "0111"; -- 0x00b
	when "000001100" => qq <= "1101"; -- 0x00c
	when "000001101" => qq <= "0111"; -- 0x00d
	when "000001110" => qq <= "0000"; -- 0x00e
	when "000001111" => qq <= "0000"; -- 0x00f
	when "000010000" => qq <= "0000"; -- 0x010
	when "000010001" => qq <= "0000"; -- 0x011
	when "000010010" => qq <= "1000"; -- 0x012
	when "000010011" => qq <= "0000"; -- 0x013
	when "000010100" => qq <= "1000"; -- 0x014
	when "000010101" => qq <= "0111"; -- 0x015
	when "000010110" => qq <= "1100"; -- 0x016
	when "000010111" => qq <= "0111"; -- 0x017
	when "000011000" => qq <= "1100"; -- 0x018
	when "000011001" => qq <= "0000"; -- 0x019
	when "000011010" => qq <= "1110"; -- 0x01a
	when "000011011" => qq <= "0011"; -- 0x01b
	when "000011100" => qq <= "1110"; -- 0x01c
	when "000011101" => qq <= "0011"; -- 0x01d
	when "000011110" => qq <= "0000"; -- 0x01e
	when "000011111" => qq <= "0000"; -- 0x01f
	when "000100000" => qq <= "0000"; -- 0x020
	when "000100001" => qq <= "0000"; -- 0x021
	when "000100010" => qq <= "0000"; -- 0x022
	when "000100011" => qq <= "0000"; -- 0x023
	when "000100100" => qq <= "1001"; -- 0x024
	when "000100101" => qq <= "0000"; -- 0x025
	when "000100110" => qq <= "1100"; -- 0x026
	when "000100111" => qq <= "1110"; -- 0x027
	when "000101000" => qq <= "1100"; -- 0x028
	when "000101001" => qq <= "0111"; -- 0x029
	when "000101010" => qq <= "1110"; -- 0x02a
	when "000101011" => qq <= "0000"; -- 0x02b
	when "000101100" => qq <= "1110"; -- 0x02c
	when "000101101" => qq <= "0011"; -- 0x02d
	when "000101110" => qq <= "0000"; -- 0x02e
	when "000101111" => qq <= "0001"; -- 0x02f
	when "000110000" => qq <= "0111"; -- 0x030
	when "000110001" => qq <= "0001"; -- 0x031
	when "000110010" => qq <= "0011"; -- 0x032
	when "000110011" => qq <= "0001"; -- 0x033
	when "000110100" => qq <= "1000"; -- 0x034
	when "000110101" => qq <= "0000"; -- 0x035
	when "000110110" => qq <= "1100"; -- 0x036
	when "000110111" => qq <= "1110"; -- 0x037
	when "000111000" => qq <= "1110"; -- 0x038
	when "000111001" => qq <= "0111"; -- 0x039
	when "000111010" => qq <= "1111"; -- 0x03a
	when "000111011" => qq <= "0000"; -- 0x03b
	when "000111100" => qq <= "1110"; -- 0x03c
	when "000111101" => qq <= "0011"; -- 0x03d
	when "000111110" => qq <= "0000"; -- 0x03e
	when "000111111" => qq <= "0001"; -- 0x03f
	when "001000000" => qq <= "1110"; -- 0x040
	when "001000001" => qq <= "1111"; -- 0x041
	when "001000010" => qq <= "0111"; -- 0x042
	when "001000011" => qq <= "0111"; -- 0x043
	when "001000100" => qq <= "0000"; -- 0x044
	when "001000101" => qq <= "0001"; -- 0x045
	when "001000110" => qq <= "1100"; -- 0x046
	when "001000111" => qq <= "1100"; -- 0x047
	when "001001000" => qq <= "1111"; -- 0x048
	when "001001001" => qq <= "1110"; -- 0x049
	when "001001010" => qq <= "1111"; -- 0x04a
	when "001001011" => qq <= "0000"; -- 0x04b
	when "001001100" => qq <= "0111"; -- 0x04c
	when "001001101" => qq <= "0001"; -- 0x04d
	when "001001110" => qq <= "0000"; -- 0x04e
	when "001001111" => qq <= "0000"; -- 0x04f
	when "001010000" => qq <= "1100"; -- 0x050
	when "001010001" => qq <= "0000"; -- 0x051
	when "001010010" => qq <= "0111"; -- 0x052
	when "001010011" => qq <= "1111"; -- 0x053
	when "001010100" => qq <= "0000"; -- 0x054
	when "001010101" => qq <= "0111"; -- 0x055
	when "001010110" => qq <= "1100"; -- 0x056
	when "001010111" => qq <= "0001"; -- 0x057
	when "001011000" => qq <= "1111"; -- 0x058
	when "001011001" => qq <= "1100"; -- 0x059
	when "001011010" => qq <= "1111"; -- 0x05a
	when "001011011" => qq <= "0111"; -- 0x05b
	when "001011100" => qq <= "0011"; -- 0x05c
	when "001011101" => qq <= "0000"; -- 0x05d
	when "001011110" => qq <= "1000"; -- 0x05e
	when "001011111" => qq <= "0000"; -- 0x05f
	when "001100000" => qq <= "1000"; -- 0x060
	when "001100001" => qq <= "0000"; -- 0x061
	when "001100010" => qq <= "1101"; -- 0x062
	when "001100011" => qq <= "0000"; -- 0x063
	when "001100100" => qq <= "0000"; -- 0x064
	when "001100101" => qq <= "1111"; -- 0x065
	when "001100110" => qq <= "1110"; -- 0x066
	when "001100111" => qq <= "0011"; -- 0x067
	when "001101000" => qq <= "1111"; -- 0x068
	when "001101001" => qq <= "0000"; -- 0x069
	when "001101010" => qq <= "0111"; -- 0x06a
	when "001101011" => qq <= "1111"; -- 0x06b
	when "001101100" => qq <= "1110"; -- 0x06c
	when "001101101" => qq <= "0111"; -- 0x06d
	when "001101110" => qq <= "1111"; -- 0x06e
	when "001101111" => qq <= "0000"; -- 0x06f
	when "001110000" => qq <= "1001"; -- 0x070
	when "001110001" => qq <= "0000"; -- 0x071
	when "001110010" => qq <= "1001"; -- 0x072
	when "001110011" => qq <= "0000"; -- 0x073
	when "001110100" => qq <= "0000"; -- 0x074
	when "001110101" => qq <= "0000"; -- 0x075
	when "001110110" => qq <= "1111"; -- 0x076
	when "001110111" => qq <= "1111"; -- 0x077
	when "001111000" => qq <= "1111"; -- 0x078
	when "001111001" => qq <= "0011"; -- 0x079
	when "001111010" => qq <= "0011"; -- 0x07a
	when "001111011" => qq <= "0000"; -- 0x07b
	when "001111100" => qq <= "0111"; -- 0x07c
	when "001111101" => qq <= "0001"; -- 0x07d
	when "001111110" => qq <= "0111"; -- 0x07e
	when "001111111" => qq <= "0001"; -- 0x07f
	when "010000000" => qq <= "0011"; -- 0x080
	when "010000001" => qq <= "0001"; -- 0x081
	when "010000010" => qq <= "0011"; -- 0x082
	when "010000011" => qq <= "0001"; -- 0x083
	when "010000100" => qq <= "0001"; -- 0x084
	when "010000101" => qq <= "0000"; -- 0x085
	when "010000110" => qq <= "1111"; -- 0x086
	when "010000111" => qq <= "1111"; -- 0x087
	when "010001000" => qq <= "1111"; -- 0x088
	when "010001001" => qq <= "1111"; -- 0x089
	when "010001010" => qq <= "0001"; -- 0x08a
	when "010001011" => qq <= "0000"; -- 0x08b
	when "010001100" => qq <= "0011"; -- 0x08c
	when "010001101" => qq <= "0001"; -- 0x08d
	when "010001110" => qq <= "0011"; -- 0x08e
	when "010001111" => qq <= "0001"; -- 0x08f
	when "010010000" => qq <= "0111"; -- 0x090
	when "010010001" => qq <= "0001"; -- 0x091
	when "010010010" => qq <= "0111"; -- 0x092
	when "010010011" => qq <= "0001"; -- 0x093
	when "010010100" => qq <= "0011"; -- 0x094
	when "010010101" => qq <= "0000"; -- 0x095
	when "010010110" => qq <= "1111"; -- 0x096
	when "010010111" => qq <= "0011"; -- 0x097
	when "010011000" => qq <= "1111"; -- 0x098
	when "010011001" => qq <= "1111"; -- 0x099
	when "010011010" => qq <= "0000"; -- 0x09a
	when "010011011" => qq <= "0000"; -- 0x09b
	when "010011100" => qq <= "1001"; -- 0x09c
	when "010011101" => qq <= "0000"; -- 0x09d
	when "010011110" => qq <= "1001"; -- 0x09e
	when "010011111" => qq <= "0000"; -- 0x09f
	when "010100000" => qq <= "1111"; -- 0x0a0
	when "010100001" => qq <= "0000"; -- 0x0a1
	when "010100010" => qq <= "1110"; -- 0x0a2
	when "010100011" => qq <= "0111"; -- 0x0a3
	when "010100100" => qq <= "0111"; -- 0x0a4
	when "010100101" => qq <= "1111"; -- 0x0a5
	when "010100110" => qq <= "1111"; -- 0x0a6
	when "010100111" => qq <= "0000"; -- 0x0a7
	when "010101000" => qq <= "1110"; -- 0x0a8
	when "010101001" => qq <= "0011"; -- 0x0a9
	when "010101010" => qq <= "0000"; -- 0x0aa
	when "010101011" => qq <= "1111"; -- 0x0ab
	when "010101100" => qq <= "1101"; -- 0x0ac
	when "010101101" => qq <= "0000"; -- 0x0ad
	when "010101110" => qq <= "1000"; -- 0x0ae
	when "010101111" => qq <= "0000"; -- 0x0af
	when "010110000" => qq <= "1000"; -- 0x0b0
	when "010110001" => qq <= "0000"; -- 0x0b1
	when "010110010" => qq <= "0011"; -- 0x0b2
	when "010110011" => qq <= "0000"; -- 0x0b3
	when "010110100" => qq <= "1111"; -- 0x0b4
	when "010110101" => qq <= "0111"; -- 0x0b5
	when "010110110" => qq <= "1111"; -- 0x0b6
	when "010110111" => qq <= "1100"; -- 0x0b7
	when "010111000" => qq <= "1100"; -- 0x0b8
	when "010111001" => qq <= "0001"; -- 0x0b9
	when "010111010" => qq <= "0000"; -- 0x0ba
	when "010111011" => qq <= "0111"; -- 0x0bb
	when "010111100" => qq <= "0111"; -- 0x0bc
	when "010111101" => qq <= "1111"; -- 0x0bd
	when "010111110" => qq <= "1100"; -- 0x0be
	when "010111111" => qq <= "0000"; -- 0x0bf
	when "011000000" => qq <= "0000"; -- 0x0c0
	when "011000001" => qq <= "0000"; -- 0x0c1
	when "011000010" => qq <= "0111"; -- 0x0c2
	when "011000011" => qq <= "0001"; -- 0x0c3
	when "011000100" => qq <= "1111"; -- 0x0c4
	when "011000101" => qq <= "0000"; -- 0x0c5
	when "011000110" => qq <= "1111"; -- 0x0c6
	when "011000111" => qq <= "1110"; -- 0x0c7
	when "011001000" => qq <= "1100"; -- 0x0c8
	when "011001001" => qq <= "1100"; -- 0x0c9
	when "011001010" => qq <= "0000"; -- 0x0ca
	when "011001011" => qq <= "0001"; -- 0x0cb
	when "011001100" => qq <= "0111"; -- 0x0cc
	when "011001101" => qq <= "0111"; -- 0x0cd
	when "011001110" => qq <= "1110"; -- 0x0ce
	when "011001111" => qq <= "1111"; -- 0x0cf
	when "011010000" => qq <= "0000"; -- 0x0d0
	when "011010001" => qq <= "0001"; -- 0x0d1
	when "011010010" => qq <= "1110"; -- 0x0d2
	when "011010011" => qq <= "0011"; -- 0x0d3
	when "011010100" => qq <= "1111"; -- 0x0d4
	when "011010101" => qq <= "0000"; -- 0x0d5
	when "011010110" => qq <= "1110"; -- 0x0d6
	when "011010111" => qq <= "0111"; -- 0x0d7
	when "011011000" => qq <= "1100"; -- 0x0d8
	when "011011001" => qq <= "1110"; -- 0x0d9
	when "011011010" => qq <= "1000"; -- 0x0da
	when "011011011" => qq <= "0000"; -- 0x0db
	when "011011100" => qq <= "0011"; -- 0x0dc
	when "011011101" => qq <= "0001"; -- 0x0dd
	when "011011110" => qq <= "0111"; -- 0x0de
	when "011011111" => qq <= "0001"; -- 0x0df
	when "011100000" => qq <= "0000"; -- 0x0e0
	when "011100001" => qq <= "0001"; -- 0x0e1
	when "011100010" => qq <= "1110"; -- 0x0e2
	when "011100011" => qq <= "0011"; -- 0x0e3
	when "011100100" => qq <= "1110"; -- 0x0e4
	when "011100101" => qq <= "0000"; -- 0x0e5
	when "011100110" => qq <= "1100"; -- 0x0e6
	when "011100111" => qq <= "0111"; -- 0x0e7
	when "011101000" => qq <= "1100"; -- 0x0e8
	when "011101001" => qq <= "1110"; -- 0x0e9
	when "011101010" => qq <= "1001"; -- 0x0ea
	when "011101011" => qq <= "0000"; -- 0x0eb
	when "011101100" => qq <= "0000"; -- 0x0ec
	when "011101101" => qq <= "0000"; -- 0x0ed
	when "011101110" => qq <= "0000"; -- 0x0ee
	when "011101111" => qq <= "0000"; -- 0x0ef
	when "011110000" => qq <= "0000"; -- 0x0f0
	when "011110001" => qq <= "0000"; -- 0x0f1
	when "011110010" => qq <= "1110"; -- 0x0f2
	when "011110011" => qq <= "0011"; -- 0x0f3
	when "011110100" => qq <= "1110"; -- 0x0f4
	when "011110101" => qq <= "0011"; -- 0x0f5
	when "011110110" => qq <= "1100"; -- 0x0f6
	when "011110111" => qq <= "0000"; -- 0x0f7
	when "011111000" => qq <= "1100"; -- 0x0f8
	when "011111001" => qq <= "0111"; -- 0x0f9
	when "011111010" => qq <= "1000"; -- 0x0fa
	when "011111011" => qq <= "0111"; -- 0x0fb
	when "011111100" => qq <= "1000"; -- 0x0fc
	when "011111101" => qq <= "0000"; -- 0x0fd
	when "011111110" => qq <= "0000"; -- 0x0fe
	when "011111111" => qq <= "0000"; -- 0x0ff
	when "100000000" => qq <= "0000"; -- 0x100
	when "100000001" => qq <= "0000"; -- 0x101
	when "100000010" => qq <= "1101"; -- 0x102
	when "100000011" => qq <= "0111"; -- 0x103
	when "100000100" => qq <= "1101"; -- 0x104
	when "100000101" => qq <= "0111"; -- 0x105
	when "100000110" => qq <= "1100"; -- 0x106
	when "100000111" => qq <= "0000"; -- 0x107
	when "100001000" => qq <= "1101"; -- 0x108
	when "100001001" => qq <= "0111"; -- 0x109
	when "100001010" => qq <= "1101"; -- 0x10a
	when "100001011" => qq <= "0111"; -- 0x10b
	when "100001100" => qq <= "1100"; -- 0x10c
	when "100001101" => qq <= "0000"; -- 0x10d
	when "100001110" => qq <= "1000"; -- 0x10e
	when "100001111" => qq <= "0000"; -- 0x10f
	when "100010000" => qq <= "0000"; -- 0x110
	when "100010001" => qq <= "0000"; -- 0x111
	when "100010010" => qq <= "1001"; -- 0x112
	when "100010011" => qq <= "1110"; -- 0x113
	when "100010100" => qq <= "1001"; -- 0x114
	when "100010101" => qq <= "1110"; -- 0x115
	when "100010110" => qq <= "1100"; -- 0x116
	when "100010111" => qq <= "0000"; -- 0x117
	when "100011000" => qq <= "1100"; -- 0x118
	when "100011001" => qq <= "0111"; -- 0x119
	when "100011010" => qq <= "1110"; -- 0x11a
	when "100011011" => qq <= "0111"; -- 0x11b
	when "100011100" => qq <= "1110"; -- 0x11c
	when "100011101" => qq <= "0000"; -- 0x11d
	when "100011110" => qq <= "1110"; -- 0x11e
	when "100011111" => qq <= "0000"; -- 0x11f
	when "100100000" => qq <= "0011"; -- 0x120
	when "100100001" => qq <= "0000"; -- 0x121
	when "100100010" => qq <= "1001"; -- 0x122
	when "100100011" => qq <= "1110"; -- 0x123
	when "100100100" => qq <= "1100"; -- 0x124
	when "100100101" => qq <= "1111"; -- 0x125
	when "100100110" => qq <= "1100"; -- 0x126
	when "100100111" => qq <= "0000"; -- 0x127
	when "100101000" => qq <= "1110"; -- 0x128
	when "100101001" => qq <= "0111"; -- 0x129
	when "100101010" => qq <= "1110"; -- 0x12a
	when "100101011" => qq <= "0011"; -- 0x12b
	when "100101100" => qq <= "1111"; -- 0x12c
	when "100101101" => qq <= "0000"; -- 0x12d
	when "100101110" => qq <= "1111"; -- 0x12e
	when "100101111" => qq <= "0000"; -- 0x12f
	when "100110000" => qq <= "0011"; -- 0x130
	when "100110001" => qq <= "0000"; -- 0x131
	when "100110010" => qq <= "0001"; -- 0x132
	when "100110011" => qq <= "0000"; -- 0x133
	when "100110100" => qq <= "1000"; -- 0x134
	when "100110101" => qq <= "0000"; -- 0x135
	when "100110110" => qq <= "1100"; -- 0x136
	when "100110111" => qq <= "1110"; -- 0x137
	when "100111000" => qq <= "1110"; -- 0x138
	when "100111001" => qq <= "0111"; -- 0x139
	when "100111010" => qq <= "1111"; -- 0x13a
	when "100111011" => qq <= "0000"; -- 0x13b
	when "100111100" => qq <= "1111"; -- 0x13c
	when "100111101" => qq <= "0001"; -- 0x13d
	when "100111110" => qq <= "0011"; -- 0x13e
	when "100111111" => qq <= "0000"; -- 0x13f
	when "101000000" => qq <= "0111"; -- 0x140
	when "101000001" => qq <= "0000"; -- 0x141
	when "101000010" => qq <= "0011"; -- 0x142
	when "101000011" => qq <= "0000"; -- 0x143
	when "101000100" => qq <= "1000"; -- 0x144
	when "101000101" => qq <= "0001"; -- 0x145
	when "101000110" => qq <= "1110"; -- 0x146
	when "101000111" => qq <= "0000"; -- 0x147
	when "101001000" => qq <= "1111"; -- 0x148
	when "101001001" => qq <= "1110"; -- 0x149
	when "101001010" => qq <= "1111"; -- 0x14a
	when "101001011" => qq <= "0111"; -- 0x14b
	when "101001100" => qq <= "0011"; -- 0x14c
	when "101001101" => qq <= "0000"; -- 0x14d
	when "101001110" => qq <= "0000"; -- 0x14e
	when "101001111" => qq <= "0000"; -- 0x14f
	when "101010000" => qq <= "1110"; -- 0x150
	when "101010001" => qq <= "0000"; -- 0x151
	when "101010010" => qq <= "0111"; -- 0x152
	when "101010011" => qq <= "0001"; -- 0x153
	when "101010100" => qq <= "0000"; -- 0x154
	when "101010101" => qq <= "0011"; -- 0x155
	when "101010110" => qq <= "1110"; -- 0x156
	when "101010111" => qq <= "0001"; -- 0x157
	when "101011000" => qq <= "1111"; -- 0x158
	when "101011001" => qq <= "1100"; -- 0x159
	when "101011010" => qq <= "0111"; -- 0x15a
	when "101011011" => qq <= "1111"; -- 0x15b
	when "101011100" => qq <= "0000"; -- 0x15c
	when "101011101" => qq <= "0000"; -- 0x15d
	when "101011110" => qq <= "1000"; -- 0x15e
	when "101011111" => qq <= "0000"; -- 0x15f
	when "101100000" => qq <= "0000"; -- 0x160
	when "101100001" => qq <= "0000"; -- 0x161
	when "101100010" => qq <= "1001"; -- 0x162
	when "101100011" => qq <= "0000"; -- 0x163
	when "101100100" => qq <= "0000"; -- 0x164
	when "101100101" => qq <= "0011"; -- 0x165
	when "101100110" => qq <= "1110"; -- 0x166
	when "101100111" => qq <= "0111"; -- 0x167
	when "101101000" => qq <= "1111"; -- 0x168
	when "101101001" => qq <= "0000"; -- 0x169
	when "101101010" => qq <= "0011"; -- 0x16a
	when "101101011" => qq <= "1111"; -- 0x16b
	when "101101100" => qq <= "1100"; -- 0x16c
	when "101101101" => qq <= "0111"; -- 0x16d
	when "101101110" => qq <= "1110"; -- 0x16e
	when "101101111" => qq <= "0000"; -- 0x16f
	when "101110000" => qq <= "0111"; -- 0x170
	when "101110001" => qq <= "0001"; -- 0x171
	when "101110010" => qq <= "0111"; -- 0x172
	when "101110011" => qq <= "0001"; -- 0x173
	when "101110100" => qq <= "0011"; -- 0x174
	when "101110101" => qq <= "0000"; -- 0x175
	when "101110110" => qq <= "1111"; -- 0x176
	when "101110111" => qq <= "0001"; -- 0x177
	when "101111000" => qq <= "1111"; -- 0x178
	when "101111001" => qq <= "0011"; -- 0x179
	when "101111010" => qq <= "1100"; -- 0x17a
	when "101111011" => qq <= "0011"; -- 0x17b
	when "101111100" => qq <= "1110"; -- 0x17c
	when "101111101" => qq <= "0111"; -- 0x17d
	when "101111110" => qq <= "1110"; -- 0x17e
	when "101111111" => qq <= "0111"; -- 0x17f
	when "110000000" => qq <= "0111"; -- 0x180
	when "110000001" => qq <= "0011"; -- 0x181
	when "110000010" => qq <= "0111"; -- 0x182
	when "110000011" => qq <= "0011"; -- 0x183
	when "110000100" => qq <= "0011"; -- 0x184
	when "110000101" => qq <= "0001"; -- 0x185
	when "110000110" => qq <= "1111"; -- 0x186
	when "110000111" => qq <= "0011"; -- 0x187
	when "110001000" => qq <= "1111"; -- 0x188
	when "110001001" => qq <= "0011"; -- 0x189
	when "110001010" => qq <= "0011"; -- 0x18a
	when "110001011" => qq <= "0001"; -- 0x18b
	when "110001100" => qq <= "0111"; -- 0x18c
	when "110001101" => qq <= "0011"; -- 0x18d
	when "110001110" => qq <= "0111"; -- 0x18e
	when "110001111" => qq <= "0011"; -- 0x18f
	when "110010000" => qq <= "1110"; -- 0x190
	when "110010001" => qq <= "0111"; -- 0x191
	when "110010010" => qq <= "1110"; -- 0x192
	when "110010011" => qq <= "0111"; -- 0x193
	when "110010100" => qq <= "1100"; -- 0x194
	when "110010101" => qq <= "0011"; -- 0x195
	when "110010110" => qq <= "1111"; -- 0x196
	when "110010111" => qq <= "0011"; -- 0x197
	when "110011000" => qq <= "1111"; -- 0x198
	when "110011001" => qq <= "0001"; -- 0x199
	when "110011010" => qq <= "0011"; -- 0x19a
	when "110011011" => qq <= "0000"; -- 0x19b
	when "110011100" => qq <= "0111"; -- 0x19c
	when "110011101" => qq <= "0001"; -- 0x19d
	when "110011110" => qq <= "0111"; -- 0x19e
	when "110011111" => qq <= "0001"; -- 0x19f
	when "110100000" => qq <= "1110"; -- 0x1a0
	when "110100001" => qq <= "0000"; -- 0x1a1
	when "110100010" => qq <= "1100"; -- 0x1a2
	when "110100011" => qq <= "0111"; -- 0x1a3
	when "110100100" => qq <= "0011"; -- 0x1a4
	when "110100101" => qq <= "1111"; -- 0x1a5
	when "110100110" => qq <= "1111"; -- 0x1a6
	when "110100111" => qq <= "0000"; -- 0x1a7
	when "110101000" => qq <= "1110"; -- 0x1a8
	when "110101001" => qq <= "0111"; -- 0x1a9
	when "110101010" => qq <= "0000"; -- 0x1aa
	when "110101011" => qq <= "0011"; -- 0x1ab
	when "110101100" => qq <= "1001"; -- 0x1ac
	when "110101101" => qq <= "0000"; -- 0x1ad
	when "110101110" => qq <= "0000"; -- 0x1ae
	when "110101111" => qq <= "0000"; -- 0x1af
	when "110110000" => qq <= "1000"; -- 0x1b0
	when "110110001" => qq <= "0000"; -- 0x1b1
	when "110110010" => qq <= "0000"; -- 0x1b2
	when "110110011" => qq <= "0000"; -- 0x1b3
	when "110110100" => qq <= "0111"; -- 0x1b4
	when "110110101" => qq <= "1111"; -- 0x1b5
	when "110110110" => qq <= "1111"; -- 0x1b6
	when "110110111" => qq <= "1100"; -- 0x1b7
	when "110111000" => qq <= "1110"; -- 0x1b8
	when "110111001" => qq <= "0001"; -- 0x1b9
	when "110111010" => qq <= "0000"; -- 0x1ba
	when "110111011" => qq <= "0011"; -- 0x1bb
	when "110111100" => qq <= "0111"; -- 0x1bc
	when "110111101" => qq <= "0001"; -- 0x1bd
	when "110111110" => qq <= "1110"; -- 0x1be
	when "110111111" => qq <= "0000"; -- 0x1bf
	when "111000000" => qq <= "0000"; -- 0x1c0
	when "111000001" => qq <= "0000"; -- 0x1c1
	when "111000010" => qq <= "0011"; -- 0x1c2
	when "111000011" => qq <= "0000"; -- 0x1c3
	when "111000100" => qq <= "1111"; -- 0x1c4
	when "111000101" => qq <= "0111"; -- 0x1c5
	when "111000110" => qq <= "1111"; -- 0x1c6
	when "111000111" => qq <= "1110"; -- 0x1c7
	when "111001000" => qq <= "1110"; -- 0x1c8
	when "111001001" => qq <= "0000"; -- 0x1c9
	when "111001010" => qq <= "1000"; -- 0x1ca
	when "111001011" => qq <= "0001"; -- 0x1cb
	when "111001100" => qq <= "0011"; -- 0x1cc
	when "111001101" => qq <= "0000"; -- 0x1cd
	when "111001110" => qq <= "0111"; -- 0x1ce
	when "111001111" => qq <= "0000"; -- 0x1cf
	when "111010000" => qq <= "0011"; -- 0x1d0
	when "111010001" => qq <= "0000"; -- 0x1d1
	when "111010010" => qq <= "1111"; -- 0x1d2
	when "111010011" => qq <= "0001"; -- 0x1d3
	when "111010100" => qq <= "1111"; -- 0x1d4
	when "111010101" => qq <= "0000"; -- 0x1d5
	when "111010110" => qq <= "1111"; -- 0x1d6
	when "111010111" => qq <= "0111"; -- 0x1d7
	when "111011000" => qq <= "1100"; -- 0x1d8
	when "111011001" => qq <= "1110"; -- 0x1d9
	when "111011010" => qq <= "1000"; -- 0x1da
	when "111011011" => qq <= "0000"; -- 0x1db
	when "111011100" => qq <= "0001"; -- 0x1dc
	when "111011101" => qq <= "0000"; -- 0x1dd
	when "111011110" => qq <= "0011"; -- 0x1de
	when "111011111" => qq <= "0000"; -- 0x1df
	when "111100000" => qq <= "0111"; -- 0x1e0
	when "111100001" => qq <= "0000"; -- 0x1e1
	when "111100010" => qq <= "1111"; -- 0x1e2
	when "111100011" => qq <= "0000"; -- 0x1e3
	when "111100100" => qq <= "1110"; -- 0x1e4
	when "111100101" => qq <= "0011"; -- 0x1e5
	when "111100110" => qq <= "1110"; -- 0x1e6
	when "111100111" => qq <= "0111"; -- 0x1e7
	when "111101000" => qq <= "1100"; -- 0x1e8
	when "111101001" => qq <= "0000"; -- 0x1e9
	when "111101010" => qq <= "1100"; -- 0x1ea
	when "111101011" => qq <= "1111"; -- 0x1eb
	when "111101100" => qq <= "1001"; -- 0x1ec
	when "111101101" => qq <= "1110"; -- 0x1ed
	when "111101110" => qq <= "0011"; -- 0x1ee
	when "111101111" => qq <= "0000"; -- 0x1ef
	when "111110000" => qq <= "1110"; -- 0x1f0
	when "111110001" => qq <= "0000"; -- 0x1f1
	when "111110010" => qq <= "1110"; -- 0x1f2
	when "111110011" => qq <= "0000"; -- 0x1f3
	when "111110100" => qq <= "1110"; -- 0x1f4
	when "111110101" => qq <= "0111"; -- 0x1f5
	when "111110110" => qq <= "1100"; -- 0x1f6
	when "111110111" => qq <= "0111"; -- 0x1f7
	when "111111000" => qq <= "1100"; -- 0x1f8
	when "111111001" => qq <= "0000"; -- 0x1f9
	when "111111010" => qq <= "1001"; -- 0x1fa
	when "111111011" => qq <= "1110"; -- 0x1fb
	when "111111100" => qq <= "1001"; -- 0x1fc
	when "111111101" => qq <= "1110"; -- 0x1fd
	when "111111110" => qq <= "0000"; -- 0x1fe
	when "111111111" => qq <= "0000"; -- 0x1ff
	when others => qq <= "0000";
END CASE; 
END PROCESS; 
END SYN; 
