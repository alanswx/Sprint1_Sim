library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
ENTITY prog_rom3 IS
PORT
(
	address         : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
	clock           : IN STD_LOGIC  := '1';
	q               : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END prog_rom3; 
ARCHITECTURE SYN OF prog_rom3 IS	
signal qq : STD_LOGIC_VECTOR (7 DOWNTO 0);
begin
q<=qq;
PROCESS (address)
begin
CASE address IS 
	when "00000000000" => qq <= "01001000"; -- 0x000
	when "00000000001" => qq <= "10001010"; -- 0x001
	when "00000000010" => qq <= "01001000"; -- 0x002
	when "00000000011" => qq <= "11011000"; -- 0x003
	when "00000000100" => qq <= "10100101"; -- 0x004
	when "00000000101" => qq <= "00110000"; -- 0x005
	when "00000000110" => qq <= "11010000"; -- 0x006
	when "00000000111" => qq <= "00000011"; -- 0x007
	when "00000001000" => qq <= "10001101"; -- 0x008
	when "00000001001" => qq <= "00000000"; -- 0x009
	when "00000001010" => qq <= "00001111"; -- 0x00a
	when "00000001011" => qq <= "00101100"; -- 0x00b
	when "00000001100" => qq <= "00101100"; -- 0x00c
	when "00000001101" => qq <= "00001000"; -- 0x00d
	when "00000001110" => qq <= "00010000"; -- 0x00e
	when "00000001111" => qq <= "00100000"; -- 0x00f
	when "00000010000" => qq <= "10100101"; -- 0x010
	when "00000010001" => qq <= "01100001"; -- 0x011
	when "00000010010" => qq <= "11001001"; -- 0x012
	when "00000010011" => qq <= "10010010"; -- 0x013
	when "00000010100" => qq <= "11010000"; -- 0x014
	when "00000010101" => qq <= "00011110"; -- 0x015
	when "00000010110" => qq <= "10100101"; -- 0x016
	when "00000010111" => qq <= "01100000"; -- 0x017
	when "00000011000" => qq <= "11001001"; -- 0x018
	when "00000011001" => qq <= "00111111"; -- 0x019
	when "00000011010" => qq <= "11010000"; -- 0x01a
	when "00000011011" => qq <= "00011000"; -- 0x01b
	when "00000011100" => qq <= "10111010"; -- 0x01c
	when "00000011101" => qq <= "10111101"; -- 0x01d
	when "00000011110" => qq <= "00000101"; -- 0x01e
	when "00000011111" => qq <= "00000001"; -- 0x01f
	when "00000100000" => qq <= "11001001"; -- 0x020
	when "00000100001" => qq <= "00100000"; -- 0x021
	when "00000100010" => qq <= "10110000"; -- 0x022
	when "00000100011" => qq <= "00001100"; -- 0x023
	when "00000100100" => qq <= "11001001"; -- 0x024
	when "00000100101" => qq <= "01000000"; -- 0x025
	when "00000100110" => qq <= "10010000"; -- 0x026
	when "00000100111" => qq <= "00001000"; -- 0x027
	when "00000101000" => qq <= "11001001"; -- 0x028
	when "00000101001" => qq <= "00010000"; -- 0x029
	when "00000101010" => qq <= "10010000"; -- 0x02a
	when "00000101011" => qq <= "00010000"; -- 0x02b
	when "00000101100" => qq <= "11001001"; -- 0x02c
	when "00000101101" => qq <= "00011000"; -- 0x02d
	when "00000101110" => qq <= "10110000"; -- 0x02e
	when "00000101111" => qq <= "00001100"; -- 0x02f
	when "00000110000" => qq <= "01101000"; -- 0x030
	when "00000110001" => qq <= "10101010"; -- 0x031
	when "00000110010" => qq <= "01101000"; -- 0x032
	when "00000110011" => qq <= "01000000"; -- 0x033
	when "00000110100" => qq <= "10101001"; -- 0x034
	when "00000110101" => qq <= "10010010"; -- 0x035
	when "00000110110" => qq <= "10000101"; -- 0x036
	when "00000110111" => qq <= "01100001"; -- 0x037
	when "00000111000" => qq <= "10101001"; -- 0x038
	when "00000111001" => qq <= "00111111"; -- 0x039
	when "00000111010" => qq <= "10000101"; -- 0x03a
	when "00000111011" => qq <= "01100000"; -- 0x03b
	when "00000111100" => qq <= "01111000"; -- 0x03c
	when "00000111101" => qq <= "11011000"; -- 0x03d
	when "00000111110" => qq <= "10100010"; -- 0x03e
	when "00000111111" => qq <= "01111111"; -- 0x03f
	when "00001000000" => qq <= "10011010"; -- 0x040
	when "00001000001" => qq <= "10101101"; -- 0x041
	when "00001000010" => qq <= "00000000"; -- 0x042
	when "00001000011" => qq <= "00011000"; -- 0x043
	when "00001000100" => qq <= "11001001"; -- 0x044
	when "00001000101" => qq <= "10101010"; -- 0x045
	when "00001000110" => qq <= "11110000"; -- 0x046
	when "00001000111" => qq <= "00000011"; -- 0x047
	when "00001001000" => qq <= "01001100"; -- 0x048
	when "00001001001" => qq <= "01001110"; -- 0x049
	when "00001001010" => qq <= "00110000"; -- 0x04a
	when "00001001011" => qq <= "00100000"; -- 0x04b
	when "00001001100" => qq <= "00000000"; -- 0x04c
	when "00001001101" => qq <= "00011000"; -- 0x04d
	when "00001001110" => qq <= "10100010"; -- 0x04e
	when "00001001111" => qq <= "00010110"; -- 0x04f
	when "00001010000" => qq <= "00100000"; -- 0x050
	when "00001010001" => qq <= "10110111"; -- 0x051
	when "00001010010" => qq <= "00111000"; -- 0x052
	when "00001010011" => qq <= "10100010"; -- 0x053
	when "00001010100" => qq <= "00000100"; -- 0x054
	when "00001010101" => qq <= "00100000"; -- 0x055
	when "00001010110" => qq <= "10110111"; -- 0x056
	when "00001010111" => qq <= "00111000"; -- 0x057
	when "00001011000" => qq <= "10100010"; -- 0x058
	when "00001011001" => qq <= "00001100"; -- 0x059
	when "00001011010" => qq <= "00100000"; -- 0x05a
	when "00001011011" => qq <= "10110111"; -- 0x05b
	when "00001011100" => qq <= "00111000"; -- 0x05c
	when "00001011101" => qq <= "00100000"; -- 0x05d
	when "00001011110" => qq <= "00000011"; -- 0x05e
	when "00001011111" => qq <= "00110111"; -- 0x05f
	when "00001100000" => qq <= "00100000"; -- 0x060
	when "00001100001" => qq <= "01101001"; -- 0x061
	when "00001100010" => qq <= "00110000"; -- 0x062
	when "00001100011" => qq <= "00100000"; -- 0x063
	when "00001100100" => qq <= "11110111"; -- 0x064
	when "00001100101" => qq <= "00110000"; -- 0x065
	when "00001100110" => qq <= "01001100"; -- 0x066
	when "00001100111" => qq <= "01100000"; -- 0x067
	when "00001101000" => qq <= "00110000"; -- 0x068
	when "00001101001" => qq <= "10101001"; -- 0x069
	when "00001101010" => qq <= "00000000"; -- 0x06a
	when "00001101011" => qq <= "10000101"; -- 0x06b
	when "00001101100" => qq <= "00110101"; -- 0x06c
	when "00001101101" => qq <= "10000101"; -- 0x06d
	when "00001101110" => qq <= "00111000"; -- 0x06e
	when "00001101111" => qq <= "10001101"; -- 0x06f
	when "00001110000" => qq <= "00000001"; -- 0x070
	when "00001110001" => qq <= "00001100"; -- 0x071
	when "00001110010" => qq <= "00100000"; -- 0x072
	when "00001110011" => qq <= "11001101"; -- 0x073
	when "00001110100" => qq <= "00111000"; -- 0x074
	when "00001110101" => qq <= "00100000"; -- 0x075
	when "00001110110" => qq <= "11011010"; -- 0x076
	when "00001110111" => qq <= "00110101"; -- 0x077
	when "00001111000" => qq <= "00100000"; -- 0x078
	when "00001111001" => qq <= "11101110"; -- 0x079
	when "00001111010" => qq <= "00111001"; -- 0x07a
	when "00001111011" => qq <= "00100000"; -- 0x07b
	when "00001111100" => qq <= "11111111"; -- 0x07c
	when "00001111101" => qq <= "00110111"; -- 0x07d
	when "00001111110" => qq <= "10101001"; -- 0x07e
	when "00001111111" => qq <= "00000001"; -- 0x07f
	when "00010000000" => qq <= "10100010"; -- 0x080
	when "00010000001" => qq <= "00011110"; -- 0x081
	when "00010000010" => qq <= "00100000"; -- 0x082
	when "00010000011" => qq <= "10001010"; -- 0x083
	when "00010000100" => qq <= "00111000"; -- 0x084
	when "00010000101" => qq <= "10101001"; -- 0x085
	when "00010000110" => qq <= "00000000"; -- 0x086
	when "00010000111" => qq <= "10100110"; -- 0x087
	when "00010001000" => qq <= "01010001"; -- 0x088
	when "00010001001" => qq <= "00100000"; -- 0x089
	when "00010001010" => qq <= "10001010"; -- 0x08a
	when "00010001011" => qq <= "00111000"; -- 0x08b
	when "00010001100" => qq <= "10101001"; -- 0x08c
	when "00010001101" => qq <= "00000000"; -- 0x08d
	when "00010001110" => qq <= "10100010"; -- 0x08e
	when "00010001111" => qq <= "00001110"; -- 0x08f
	when "00010010000" => qq <= "00100000"; -- 0x090
	when "00010010001" => qq <= "10001010"; -- 0x091
	when "00010010010" => qq <= "00111000"; -- 0x092
	when "00010010011" => qq <= "10101001"; -- 0x093
	when "00010010100" => qq <= "00000000"; -- 0x094
	when "00010010101" => qq <= "10100010"; -- 0x095
	when "00010010110" => qq <= "00010000"; -- 0x096
	when "00010010111" => qq <= "00100000"; -- 0x097
	when "00010011000" => qq <= "10001010"; -- 0x098
	when "00010011001" => qq <= "00111000"; -- 0x099
	when "00010011010" => qq <= "11100110"; -- 0x09a
	when "00010011011" => qq <= "00110000"; -- 0x09b
	when "00010011100" => qq <= "10101101"; -- 0x09c
	when "00010011101" => qq <= "00110000"; -- 0x09d
	when "00010011110" => qq <= "00000000"; -- 0x09e
	when "00010011111" => qq <= "11010000"; -- 0x09f
	when "00010100000" => qq <= "00010001"; -- 0x0a0
	when "00010100001" => qq <= "11100110"; -- 0x0a1
	when "00010100010" => qq <= "00110101"; -- 0x0a2
	when "00010100011" => qq <= "10100101"; -- 0x0a3
	when "00010100100" => qq <= "00110101"; -- 0x0a4
	when "00010100101" => qq <= "11001001"; -- 0x0a5
	when "00010100110" => qq <= "00001100"; -- 0x0a6
	when "00010100111" => qq <= "11010000"; -- 0x0a7
	when "00010101000" => qq <= "00001001"; -- 0x0a8
	when "00010101001" => qq <= "10101001"; -- 0x0a9
	when "00010101010" => qq <= "00000000"; -- 0x0aa
	when "00010101011" => qq <= "10000101"; -- 0x0ab
	when "00010101100" => qq <= "00110101"; -- 0x0ac
	when "00010101101" => qq <= "10000101"; -- 0x0ad
	when "00010101110" => qq <= "00111000"; -- 0x0ae
	when "00010101111" => qq <= "01001100"; -- 0x0af
	when "00010110000" => qq <= "01110010"; -- 0x0b0
	when "00010110001" => qq <= "00110000"; -- 0x0b1
	when "00010110010" => qq <= "00101100"; -- 0x0b2
	when "00010110011" => qq <= "00101100"; -- 0x0b3
	when "00010110100" => qq <= "00001000"; -- 0x0b4
	when "00010110101" => qq <= "00110000"; -- 0x0b5
	when "00010110110" => qq <= "00000011"; -- 0x0b6
	when "00010110111" => qq <= "01001100"; -- 0x0b7
	when "00010111000" => qq <= "01010010"; -- 0x0b8
	when "00010111001" => qq <= "00111010"; -- 0x0b9
	when "00010111010" => qq <= "00100000"; -- 0x0ba
	when "00010111011" => qq <= "00111101"; -- 0x0bb
	when "00010111100" => qq <= "00111010"; -- 0x0bc
	when "00010111101" => qq <= "10100010"; -- 0x0bd
	when "00010111110" => qq <= "00000000"; -- 0x0be
	when "00010111111" => qq <= "00100000"; -- 0x0bf
	when "00011000000" => qq <= "10000101"; -- 0x0c0
	when "00011000001" => qq <= "00110100"; -- 0x0c1
	when "00011000010" => qq <= "11101000"; -- 0x0c2
	when "00011000011" => qq <= "11100000"; -- 0x0c3
	when "00011000100" => qq <= "00000100"; -- 0x0c4
	when "00011000101" => qq <= "11010000"; -- 0x0c5
	when "00011000110" => qq <= "11111000"; -- 0x0c6
	when "00011000111" => qq <= "10101001"; -- 0x0c7
	when "00011001000" => qq <= "00000000"; -- 0x0c8
	when "00011001001" => qq <= "10000101"; -- 0x0c9
	when "00011001010" => qq <= "00010110"; -- 0x0ca
	when "00011001011" => qq <= "10001101"; -- 0x0cb
	when "00011001100" => qq <= "00010100"; -- 0x0cc
	when "00011001101" => qq <= "00000000"; -- 0x0cd
	when "00011001110" => qq <= "10001101"; -- 0x0ce
	when "00011001111" => qq <= "00010000"; -- 0x0cf
	when "00011010000" => qq <= "00001100"; -- 0x0d0
	when "00011010001" => qq <= "00101100"; -- 0x0d1
	when "00011010010" => qq <= "01000000"; -- 0x0d2
	when "00011010011" => qq <= "00001000"; -- 0x0d3
	when "00011010100" => qq <= "00010000"; -- 0x0d4
	when "00011010101" => qq <= "00000010"; -- 0x0d5
	when "00011010110" => qq <= "01110000"; -- 0x0d6
	when "00011010111" => qq <= "00000011"; -- 0x0d7
	when "00011011000" => qq <= "00100000"; -- 0x0d8
	when "00011011001" => qq <= "11111111"; -- 0x0d9
	when "00011011010" => qq <= "00110111"; -- 0x0da
	when "00011011011" => qq <= "00101100"; -- 0x0db
	when "00011011100" => qq <= "00000000"; -- 0x0dc
	when "00011011101" => qq <= "00001100"; -- 0x0dd
	when "00011011110" => qq <= "01010000"; -- 0x0de
	when "00011011111" => qq <= "11110001"; -- 0x0df
	when "00011100000" => qq <= "10001101"; -- 0x0e0
	when "00011100001" => qq <= "10000000"; -- 0x0e1
	when "00011100010" => qq <= "00001100"; -- 0x0e2
	when "00011100011" => qq <= "10100101"; -- 0x0e3
	when "00011100100" => qq <= "00110110"; -- 0x0e4
	when "00011100101" => qq <= "11010000"; -- 0x0e5
	when "00011100110" => qq <= "00000100"; -- 0x0e6
	when "00011100111" => qq <= "10100101"; -- 0x0e7
	when "00011101000" => qq <= "00100000"; -- 0x0e8
	when "00011101001" => qq <= "11110000"; -- 0x0e9
	when "00011101010" => qq <= "10101111"; -- 0x0ea
	when "00011101011" => qq <= "00100000"; -- 0x0eb
	when "00011101100" => qq <= "10111010"; -- 0x0ec
	when "00011101101" => qq <= "00111001"; -- 0x0ed
	when "00011101110" => qq <= "10100101"; -- 0x0ee
	when "00011101111" => qq <= "00110110"; -- 0x0ef
	when "00011110000" => qq <= "11010000"; -- 0x0f0
	when "00011110001" => qq <= "00000100"; -- 0x0f1
	when "00011110010" => qq <= "10100101"; -- 0x0f2
	when "00011110011" => qq <= "00100000"; -- 0x0f3
	when "00011110100" => qq <= "11110000"; -- 0x0f4
	when "00011110101" => qq <= "10100100"; -- 0x0f5
	when "00011110110" => qq <= "01100000"; -- 0x0f6
	when "00011110111" => qq <= "11101010"; -- 0x0f7
	when "00011111000" => qq <= "10100010"; -- 0x0f8
	when "00011111001" => qq <= "00000000"; -- 0x0f9
	when "00011111010" => qq <= "10000110"; -- 0x0fa
	when "00011111011" => qq <= "00110101"; -- 0x0fb
	when "00011111100" => qq <= "10000110"; -- 0x0fc
	when "00011111101" => qq <= "00111000"; -- 0x0fd
	when "00011111110" => qq <= "00100000"; -- 0x0fe
	when "00011111111" => qq <= "11001101"; -- 0x0ff
	when "00100000000" => qq <= "00111000"; -- 0x100
	when "00100000001" => qq <= "10100010"; -- 0x101
	when "00100000010" => qq <= "00000110"; -- 0x102
	when "00100000011" => qq <= "00100000"; -- 0x103
	when "00100000100" => qq <= "10110111"; -- 0x104
	when "00100000101" => qq <= "00111000"; -- 0x105
	when "00100000110" => qq <= "10101001"; -- 0x106
	when "00100000111" => qq <= "00000000"; -- 0x107
	when "00100001000" => qq <= "10100010"; -- 0x108
	when "00100001001" => qq <= "00000000"; -- 0x109
	when "00100001010" => qq <= "00100000"; -- 0x10a
	when "00100001011" => qq <= "10001010"; -- 0x10b
	when "00100001100" => qq <= "00111000"; -- 0x10c
	when "00100001101" => qq <= "10101001"; -- 0x10d
	when "00100001110" => qq <= "00000000"; -- 0x10e
	when "00100001111" => qq <= "10000101"; -- 0x10f
	when "00100010000" => qq <= "00101010"; -- 0x110
	when "00100010001" => qq <= "00100000"; -- 0x111
	when "00100010010" => qq <= "11011010"; -- 0x112
	when "00100010011" => qq <= "00110101"; -- 0x113
	when "00100010100" => qq <= "00100000"; -- 0x114
	when "00100010101" => qq <= "00111101"; -- 0x115
	when "00100010110" => qq <= "00111010"; -- 0x116
	when "00100010111" => qq <= "00100000"; -- 0x117
	when "00100011000" => qq <= "11111111"; -- 0x118
	when "00100011001" => qq <= "00110111"; -- 0x119
	when "00100011010" => qq <= "10001101"; -- 0x11a
	when "00100011011" => qq <= "10000000"; -- 0x11b
	when "00100011100" => qq <= "00001100"; -- 0x11c
	when "00100011101" => qq <= "10100101"; -- 0x11d
	when "00100011110" => qq <= "00100000"; -- 0x11e
	when "00100011111" => qq <= "11110000"; -- 0x11f
	when "00100100000" => qq <= "11110110"; -- 0x120
	when "00100100001" => qq <= "10001101"; -- 0x121
	when "00100100010" => qq <= "00110001"; -- 0x122
	when "00100100011" => qq <= "00001100"; -- 0x123
	when "00100100100" => qq <= "10101001"; -- 0x124
	when "00100100101" => qq <= "00000000"; -- 0x125
	when "00100100110" => qq <= "10100010"; -- 0x126
	when "00100100111" => qq <= "00010100"; -- 0x127
	when "00100101000" => qq <= "00100000"; -- 0x128
	when "00100101001" => qq <= "10001010"; -- 0x129
	when "00100101010" => qq <= "00111000"; -- 0x12a
	when "00100101011" => qq <= "00101100"; -- 0x12b
	when "00100101100" => qq <= "00101101"; -- 0x12c
	when "00100101101" => qq <= "00001000"; -- 0x12d
	when "00100101110" => qq <= "00110000"; -- 0x12e
	when "00100101111" => qq <= "11100111"; -- 0x12f
	when "00100110000" => qq <= "11000110"; -- 0x130
	when "00100110001" => qq <= "00100000"; -- 0x131
	when "00100110010" => qq <= "10100010"; -- 0x132
	when "00100110011" => qq <= "00000000"; -- 0x133
	when "00100110100" => qq <= "00100000"; -- 0x134
	when "00100110101" => qq <= "10110111"; -- 0x135
	when "00100110110" => qq <= "00111000"; -- 0x136
	when "00100110111" => qq <= "10100010"; -- 0x137
	when "00100111000" => qq <= "00010100"; -- 0x138
	when "00100111001" => qq <= "00100000"; -- 0x139
	when "00100111010" => qq <= "10110111"; -- 0x13a
	when "00100111011" => qq <= "00111000"; -- 0x13b
	when "00100111100" => qq <= "10100010"; -- 0x13c
	when "00100111101" => qq <= "00010010"; -- 0x13d
	when "00100111110" => qq <= "00100000"; -- 0x13e
	when "00100111111" => qq <= "10110111"; -- 0x13f
	when "00101000000" => qq <= "00111000"; -- 0x140
	when "00101000001" => qq <= "10100101"; -- 0x141
	when "00101000010" => qq <= "00111010"; -- 0x142
	when "00101000011" => qq <= "11001001"; -- 0x143
	when "00101000100" => qq <= "01000000"; -- 0x144
	when "00101000101" => qq <= "11110000"; -- 0x145
	when "00101000110" => qq <= "00010101"; -- 0x146
	when "00101000111" => qq <= "10101001"; -- 0x147
	when "00101001000" => qq <= "00000000"; -- 0x148
	when "00101001001" => qq <= "10100010"; -- 0x149
	when "00101001010" => qq <= "00010010"; -- 0x14a
	when "00101001011" => qq <= "00100000"; -- 0x14b
	when "00101001100" => qq <= "10001010"; -- 0x14c
	when "00101001101" => qq <= "00111000"; -- 0x14d
	when "00101001110" => qq <= "10100101"; -- 0x14e
	when "00101001111" => qq <= "00111010"; -- 0x14f
	when "00101010000" => qq <= "11001001"; -- 0x150
	when "00101010001" => qq <= "00110000"; -- 0x151
	when "00101010010" => qq <= "11110000"; -- 0x152
	when "00101010011" => qq <= "00000011"; -- 0x153
	when "00101010100" => qq <= "10001101"; -- 0x154
	when "00101010101" => qq <= "01110100"; -- 0x155
	when "00101010110" => qq <= "00000111"; -- 0x156
	when "00101010111" => qq <= "10100101"; -- 0x157
	when "00101011000" => qq <= "00111011"; -- 0x158
	when "00101011001" => qq <= "10001101"; -- 0x159
	when "00101011010" => qq <= "01110101"; -- 0x15a
	when "00101011011" => qq <= "00000111"; -- 0x15b
	when "00101011100" => qq <= "10001101"; -- 0x15c
	when "00101011101" => qq <= "00000000"; -- 0x15d
	when "00101011110" => qq <= "00001100"; -- 0x15e
	when "00101011111" => qq <= "00100000"; -- 0x15f
	when "00101100000" => qq <= "00111101"; -- 0x160
	when "00101100001" => qq <= "00111010"; -- 0x161
	when "00101100010" => qq <= "10100101"; -- 0x162
	when "00101100011" => qq <= "00111000"; -- 0x163
	when "00101100100" => qq <= "11110000"; -- 0x164
	when "00101100101" => qq <= "00000011"; -- 0x165
	when "00101100110" => qq <= "00100000"; -- 0x166
	when "00101100111" => qq <= "11001101"; -- 0x167
	when "00101101000" => qq <= "00111000"; -- 0x168
	when "00101101001" => qq <= "11100110"; -- 0x169
	when "00101101010" => qq <= "00110000"; -- 0x16a
	when "00101101011" => qq <= "00100000"; -- 0x16b
	when "00101101100" => qq <= "11011000"; -- 0x16c
	when "00101101101" => qq <= "00110111"; -- 0x16d
	when "00101101110" => qq <= "10100010"; -- 0x16e
	when "00101101111" => qq <= "00000001"; -- 0x16f
	when "00101110000" => qq <= "00100000"; -- 0x170
	when "00101110001" => qq <= "10000101"; -- 0x171
	when "00101110010" => qq <= "00110100"; -- 0x172
	when "00101110011" => qq <= "11101000"; -- 0x173
	when "00101110100" => qq <= "11100000"; -- 0x174
	when "00101110101" => qq <= "00000100"; -- 0x175
	when "00101110110" => qq <= "11010000"; -- 0x176
	when "00101110111" => qq <= "11111000"; -- 0x177
	when "00101111000" => qq <= "10001101"; -- 0x178
	when "00101111001" => qq <= "00010000"; -- 0x179
	when "00101111010" => qq <= "00001100"; -- 0x17a
	when "00101111011" => qq <= "10100010"; -- 0x17b
	when "00101111100" => qq <= "00000000"; -- 0x17c
	when "00101111101" => qq <= "00101100"; -- 0x17d
	when "00101111110" => qq <= "00000000"; -- 0x17e
	when "00101111111" => qq <= "00010000"; -- 0x17f
	when "00110000000" => qq <= "00110000"; -- 0x180
	when "00110000001" => qq <= "00001001"; -- 0x181
	when "00110000010" => qq <= "10100101"; -- 0x182
	when "00110000011" => qq <= "00111101"; -- 0x183
	when "00110000100" => qq <= "11110000"; -- 0x184
	when "00110000101" => qq <= "00000101"; -- 0x185
	when "00110000110" => qq <= "11000110"; -- 0x186
	when "00110000111" => qq <= "00111101"; -- 0x187
	when "00110001000" => qq <= "01001100"; -- 0x188
	when "00110001001" => qq <= "10101111"; -- 0x189
	when "00110001010" => qq <= "00110001"; -- 0x18a
	when "00110001011" => qq <= "00101100"; -- 0x18b
	when "00110001100" => qq <= "00000000"; -- 0x18c
	when "00110001101" => qq <= "00010000"; -- 0x18d
	when "00110001110" => qq <= "00110000"; -- 0x18e
	when "00110001111" => qq <= "00001001"; -- 0x18f
	when "00110010000" => qq <= "10101001"; -- 0x190
	when "00110010001" => qq <= "00000000"; -- 0x191
	when "00110010010" => qq <= "10000101"; -- 0x192
	when "00110010011" => qq <= "00111101"; -- 0x193
	when "00110010100" => qq <= "10000101"; -- 0x194
	when "00110010101" => qq <= "00111110"; -- 0x195
	when "00110010110" => qq <= "01001100"; -- 0x196
	when "00110010111" => qq <= "10101111"; -- 0x197
	when "00110011000" => qq <= "00110001"; -- 0x198
	when "00110011001" => qq <= "10101001"; -- 0x199
	when "00110011010" => qq <= "00000000"; -- 0x19a
	when "00110011011" => qq <= "10000101"; -- 0x19b
	when "00110011100" => qq <= "00110011"; -- 0x19c
	when "00110011101" => qq <= "10100101"; -- 0x19d
	when "00110011110" => qq <= "00111110"; -- 0x19e
	when "00110011111" => qq <= "11010000"; -- 0x19f
	when "00110100000" => qq <= "00001010"; -- 0x1a0
	when "00110100001" => qq <= "10101001"; -- 0x1a1
	when "00110100010" => qq <= "00000001"; -- 0x1a2
	when "00110100011" => qq <= "10010101"; -- 0x1a3
	when "00110100100" => qq <= "00000000"; -- 0x1a4
	when "00110100101" => qq <= "10000101"; -- 0x1a5
	when "00110100110" => qq <= "00111110"; -- 0x1a6
	when "00110100111" => qq <= "10101001"; -- 0x1a7
	when "00110101000" => qq <= "00001111"; -- 0x1a8
	when "00110101001" => qq <= "10000101"; -- 0x1a9
	when "00110101010" => qq <= "00010110"; -- 0x1aa
	when "00110101011" => qq <= "10101001"; -- 0x1ab
	when "00110101100" => qq <= "00010000"; -- 0x1ac
	when "00110101101" => qq <= "10000101"; -- 0x1ad
	when "00110101110" => qq <= "00111101"; -- 0x1ae
	when "00110101111" => qq <= "10100101"; -- 0x1af
	when "00110110000" => qq <= "00010110"; -- 0x1b0
	when "00110110001" => qq <= "11110000"; -- 0x1b1
	when "00110110010" => qq <= "00001010"; -- 0x1b2
	when "00110110011" => qq <= "10100101"; -- 0x1b3
	when "00110110100" => qq <= "00110000"; -- 0x1b4
	when "00110110101" => qq <= "01001010"; -- 0x1b5
	when "00110110110" => qq <= "10010000"; -- 0x1b6
	when "00110110111" => qq <= "00000101"; -- 0x1b7
	when "00110111000" => qq <= "01001010"; -- 0x1b8
	when "00110111001" => qq <= "10010000"; -- 0x1b9
	when "00110111010" => qq <= "00000010"; -- 0x1ba
	when "00110111011" => qq <= "11000110"; -- 0x1bb
	when "00110111100" => qq <= "00010110"; -- 0x1bc
	when "00110111101" => qq <= "10100101"; -- 0x1bd
	when "00110111110" => qq <= "00110011"; -- 0x1be
	when "00110111111" => qq <= "11110000"; -- 0x1bf
	when "00111000000" => qq <= "00011000"; -- 0x1c0
	when "00111000001" => qq <= "10001101"; -- 0x1c1
	when "00111000010" => qq <= "00010001"; -- 0x1c2
	when "00111000011" => qq <= "00001100"; -- 0x1c3
	when "00111000100" => qq <= "11000110"; -- 0x1c4
	when "00111000101" => qq <= "00110011"; -- 0x1c5
	when "00111000110" => qq <= "10001010"; -- 0x1c6
	when "00111000111" => qq <= "00001010"; -- 0x1c7
	when "00111001000" => qq <= "10101000"; -- 0x1c8
	when "00111001001" => qq <= "10101001"; -- 0x1c9
	when "00111001010" => qq <= "00000010"; -- 0x1ca
	when "00111001011" => qq <= "00101100"; -- 0x1cb
	when "00111001100" => qq <= "10000000"; -- 0x1cc
	when "00111001101" => qq <= "00001000"; -- 0x1cd
	when "00111001110" => qq <= "01110000"; -- 0x1ce
	when "00111001111" => qq <= "00000010"; -- 0x1cf
	when "00111010000" => qq <= "10101001"; -- 0x1d0
	when "00111010001" => qq <= "11111110"; -- 0x1d1
	when "00111010010" => qq <= "00011000"; -- 0x1d2
	when "00111010011" => qq <= "01111001"; -- 0x1d3
	when "00111010100" => qq <= "00011001"; -- 0x1d4
	when "00111010101" => qq <= "00000000"; -- 0x1d5
	when "00111010110" => qq <= "10011001"; -- 0x1d6
	when "00111010111" => qq <= "00011001"; -- 0x1d7
	when "00111011000" => qq <= "00000000"; -- 0x1d8
	when "00111011001" => qq <= "00101100"; -- 0x1d9
	when "00111011010" => qq <= "00000000"; -- 0x1da
	when "00111011011" => qq <= "00010000"; -- 0x1db
	when "00111011100" => qq <= "01010000"; -- 0x1dc
	when "00111011101" => qq <= "00000100"; -- 0x1dd
	when "00111011110" => qq <= "10101001"; -- 0x1de
	when "00111011111" => qq <= "00100000"; -- 0x1df
	when "00111100000" => qq <= "10000101"; -- 0x1e0
	when "00111100001" => qq <= "00110011"; -- 0x1e1
	when "00111100010" => qq <= "10001101"; -- 0x1e2
	when "00111100011" => qq <= "00000000"; -- 0x1e3
	when "00111100100" => qq <= "00001101"; -- 0x1e4
	when "00111100101" => qq <= "10100101"; -- 0x1e5
	when "00111100110" => qq <= "00110000"; -- 0x1e6
	when "00111100111" => qq <= "01001010"; -- 0x1e7
	when "00111101000" => qq <= "10010000"; -- 0x1e8
	when "00111101001" => qq <= "00011010"; -- 0x1e9
	when "00111101010" => qq <= "01001010"; -- 0x1ea
	when "00111101011" => qq <= "10010000"; -- 0x1eb
	when "00111101100" => qq <= "00010111"; -- 0x1ec
	when "00111101101" => qq <= "00100000"; -- 0x1ed
	when "00111101110" => qq <= "10000010"; -- 0x1ee
	when "00111101111" => qq <= "00110111"; -- 0x1ef
	when "00111110000" => qq <= "10000101"; -- 0x1f0
	when "00111110001" => qq <= "00100100"; -- 0x1f1
	when "00111110010" => qq <= "11001001"; -- 0x1f2
	when "00111110011" => qq <= "11111001"; -- 0x1f3
	when "00111110100" => qq <= "00010000"; -- 0x1f4
	when "00111110101" => qq <= "00000011"; -- 0x1f5
	when "00111110110" => qq <= "10001101"; -- 0x1f6
	when "00111110111" => qq <= "00010001"; -- 0x1f7
	when "00111111000" => qq <= "00001100"; -- 0x1f8
	when "00111111001" => qq <= "10100101"; -- 0x1f9
	when "00111111010" => qq <= "00100100"; -- 0x1fa
	when "00111111011" => qq <= "00011000"; -- 0x1fb
	when "00111111100" => qq <= "01110101"; -- 0x1fc
	when "00111111101" => qq <= "00000000"; -- 0x1fd
	when "00111111110" => qq <= "11010000"; -- 0x1fe
	when "00111111111" => qq <= "00000010"; -- 0x1ff
	when "01000000000" => qq <= "10101001"; -- 0x200
	when "01000000001" => qq <= "00000001"; -- 0x201
	when "01000000010" => qq <= "10010101"; -- 0x202
	when "01000000011" => qq <= "00000000"; -- 0x203
	when "01000000100" => qq <= "10110101"; -- 0x204
	when "01000000101" => qq <= "00000000"; -- 0x205
	when "01000000110" => qq <= "01001010"; -- 0x206
	when "01000000111" => qq <= "01001010"; -- 0x207
	when "01000001000" => qq <= "01001010"; -- 0x208
	when "01000001001" => qq <= "10000101"; -- 0x209
	when "01000001010" => qq <= "00100010"; -- 0x20a
	when "01000001011" => qq <= "10100100"; -- 0x20b
	when "01000001100" => qq <= "00110010"; -- 0x20c
	when "01000001101" => qq <= "10100101"; -- 0x20d
	when "01000001110" => qq <= "00110010"; -- 0x20e
	when "01000001111" => qq <= "00001010"; -- 0x20f
	when "01000010000" => qq <= "10000101"; -- 0x210
	when "01000010001" => qq <= "00100100"; -- 0x211
	when "01000010010" => qq <= "10111001"; -- 0x212
	when "01000010011" => qq <= "10100001"; -- 0x213
	when "01000010100" => qq <= "00111100"; -- 0x214
	when "01000010101" => qq <= "10101000"; -- 0x215
	when "01000010110" => qq <= "10101001"; -- 0x216
	when "01000010111" => qq <= "00000000"; -- 0x217
	when "01000011000" => qq <= "00011000"; -- 0x218
	when "01000011001" => qq <= "01100101"; -- 0x219
	when "01000011010" => qq <= "00100010"; -- 0x21a
	when "01000011011" => qq <= "10001000"; -- 0x21b
	when "01000011100" => qq <= "11010000"; -- 0x21c
	when "01000011101" => qq <= "11111010"; -- 0x21d
	when "01000011110" => qq <= "01001010"; -- 0x21e
	when "01000011111" => qq <= "01001010"; -- 0x21f
	when "01000100000" => qq <= "01001010"; -- 0x220
	when "01000100001" => qq <= "00111000"; -- 0x221
	when "01000100010" => qq <= "11100101"; -- 0x222
	when "01000100011" => qq <= "00100100"; -- 0x223
	when "01000100100" => qq <= "00010000"; -- 0x224
	when "01000100101" => qq <= "00000010"; -- 0x225
	when "01000100110" => qq <= "10101001"; -- 0x226
	when "01000100111" => qq <= "00000000"; -- 0x227
	when "01000101000" => qq <= "11001001"; -- 0x228
	when "01000101001" => qq <= "00010000"; -- 0x229
	when "01000101010" => qq <= "00110000"; -- 0x22a
	when "01000101011" => qq <= "00000010"; -- 0x22b
	when "01000101100" => qq <= "10101001"; -- 0x22c
	when "01000101101" => qq <= "00001111"; -- 0x22d
	when "01000101110" => qq <= "10000101"; -- 0x22e
	when "01000101111" => qq <= "00010100"; -- 0x22f
	when "01000110000" => qq <= "10001010"; -- 0x230
	when "01000110001" => qq <= "00001010"; -- 0x231
	when "01000110010" => qq <= "10101000"; -- 0x232
	when "01000110011" => qq <= "00100000"; -- 0x233
	when "01000110100" => qq <= "11011000"; -- 0x234
	when "01000110101" => qq <= "00110111"; -- 0x235
	when "01000110110" => qq <= "10110101"; -- 0x236
	when "01000110111" => qq <= "00000000"; -- 0x237
	when "01000111000" => qq <= "01001001"; -- 0x238
	when "01000111001" => qq <= "11111111"; -- 0x239
	when "01000111010" => qq <= "01001010"; -- 0x23a
	when "01000111011" => qq <= "01001010"; -- 0x23b
	when "01000111100" => qq <= "01001010"; -- 0x23c
	when "01000111101" => qq <= "01001010"; -- 0x23d
	when "01000111110" => qq <= "01001010"; -- 0x23e
	when "01000111111" => qq <= "01001010"; -- 0x23f
	when "01001000000" => qq <= "10000101"; -- 0x240
	when "01001000001" => qq <= "00100110"; -- 0x241
	when "01001000010" => qq <= "00011000"; -- 0x242
	when "01001000011" => qq <= "01101001"; -- 0x243
	when "01001000100" => qq <= "00000011"; -- 0x244
	when "01001000101" => qq <= "10000101"; -- 0x245
	when "01001000110" => qq <= "00100010"; -- 0x246
	when "01001000111" => qq <= "10111001"; -- 0x247
	when "01001001000" => qq <= "00011001"; -- 0x248
	when "01001001001" => qq <= "00000000"; -- 0x249
	when "01001001010" => qq <= "00101001"; -- 0x24a
	when "01001001011" => qq <= "11111000"; -- 0x24b
	when "01001001100" => qq <= "10000101"; -- 0x24c
	when "01001001101" => qq <= "00100100"; -- 0x24d
	when "01001001110" => qq <= "10110101"; -- 0x24e
	when "01001001111" => qq <= "00000100"; -- 0x24f
	when "01001010000" => qq <= "00101001"; -- 0x250
	when "01001010001" => qq <= "11111000"; -- 0x251
	when "01001010010" => qq <= "00111000"; -- 0x252
	when "01001010011" => qq <= "11100101"; -- 0x253
	when "01001010100" => qq <= "00100100"; -- 0x254
	when "01001010101" => qq <= "11110000"; -- 0x255
	when "01001010110" => qq <= "00100001"; -- 0x256
	when "01001010111" => qq <= "00110000"; -- 0x257
	when "01001011000" => qq <= "00010001"; -- 0x258
	when "01001011001" => qq <= "11001001"; -- 0x259
	when "01001011010" => qq <= "00010000"; -- 0x25a
	when "01001011011" => qq <= "00110000"; -- 0x25b
	when "01001011100" => qq <= "00000011"; -- 0x25c
	when "01001011101" => qq <= "10001101"; -- 0x25d
	when "01001011110" => qq <= "00010001"; -- 0x25e
	when "01001011111" => qq <= "00001100"; -- 0x25f
	when "01001100000" => qq <= "10101001"; -- 0x260
	when "01001100001" => qq <= "00000000"; -- 0x261
	when "01001100010" => qq <= "00111000"; -- 0x262
	when "01001100011" => qq <= "11100101"; -- 0x263
	when "01001100100" => qq <= "00100010"; -- 0x264
	when "01001100101" => qq <= "10000101"; -- 0x265
	when "01001100110" => qq <= "00100010"; -- 0x266
	when "01001100111" => qq <= "01001100"; -- 0x267
	when "01001101000" => qq <= "01110001"; -- 0x268
	when "01001101001" => qq <= "00110010"; -- 0x269
	when "01001101010" => qq <= "11001001"; -- 0x26a
	when "01001101011" => qq <= "11111000"; -- 0x26b
	when "01001101100" => qq <= "00010000"; -- 0x26c
	when "01001101101" => qq <= "00000011"; -- 0x26d
	when "01001101110" => qq <= "10001101"; -- 0x26e
	when "01001101111" => qq <= "00010001"; -- 0x26f
	when "01001110000" => qq <= "00001100"; -- 0x270
	when "01001110001" => qq <= "10100101"; -- 0x271
	when "01001110010" => qq <= "00100010"; -- 0x272
	when "01001110011" => qq <= "00011000"; -- 0x273
	when "01001110100" => qq <= "01110101"; -- 0x274
	when "01001110101" => qq <= "00000100"; -- 0x275
	when "01001110110" => qq <= "10010101"; -- 0x276
	when "01001110111" => qq <= "00000100"; -- 0x277
	when "01001111000" => qq <= "00100000"; -- 0x278
	when "01001111001" => qq <= "00010000"; -- 0x279
	when "01001111010" => qq <= "00110101"; -- 0x27a
	when "01001111011" => qq <= "10100101"; -- 0x27b
	when "01001111100" => qq <= "00110101"; -- 0x27c
	when "01001111101" => qq <= "00001010"; -- 0x27d
	when "01001111110" => qq <= "10101010"; -- 0x27e
	when "01001111111" => qq <= "10111101"; -- 0x27f
	when "01010000000" => qq <= "11001010"; -- 0x280
	when "01010000001" => qq <= "00101101"; -- 0x281
	when "01010000010" => qq <= "10000101"; -- 0x282
	when "01010000011" => qq <= "00100100"; -- 0x283
	when "01010000100" => qq <= "10111101"; -- 0x284
	when "01010000101" => qq <= "11001011"; -- 0x285
	when "01010000110" => qq <= "00101101"; -- 0x286
	when "01010000111" => qq <= "10000101"; -- 0x287
	when "01010001000" => qq <= "00100101"; -- 0x288
	when "01010001001" => qq <= "10101101"; -- 0x289
	when "01010001010" => qq <= "00101010"; -- 0x28a
	when "01010001011" => qq <= "00000100"; -- 0x28b
	when "01010001100" => qq <= "01001010"; -- 0x28c
	when "01010001101" => qq <= "00101001"; -- 0x28d
	when "01010001110" => qq <= "00000111"; -- 0x28e
	when "01010001111" => qq <= "00001010"; -- 0x28f
	when "01010010000" => qq <= "10101000"; -- 0x290
	when "01010010001" => qq <= "10110001"; -- 0x291
	when "01010010010" => qq <= "00100100"; -- 0x292
	when "01010010011" => qq <= "10000101"; -- 0x293
	when "01010010100" => qq <= "00101000"; -- 0x294
	when "01010010101" => qq <= "11001000"; -- 0x295
	when "01010010110" => qq <= "10110001"; -- 0x296
	when "01010010111" => qq <= "00100100"; -- 0x297
	when "01010011000" => qq <= "10000101"; -- 0x298
	when "01010011001" => qq <= "00101001"; -- 0x299
	when "01010011010" => qq <= "10100110"; -- 0x29a
	when "01010011011" => qq <= "00100010"; -- 0x29b
	when "01010011100" => qq <= "10110101"; -- 0x29c
	when "01010011101" => qq <= "01000100"; -- 0x29d
	when "01010011110" => qq <= "00101001"; -- 0x29e
	when "01010011111" => qq <= "11110000"; -- 0x29f
	when "01010100000" => qq <= "10000101"; -- 0x2a0
	when "01010100001" => qq <= "00101010"; -- 0x2a1
	when "01010100010" => qq <= "10110101"; -- 0x2a2
	when "01010100011" => qq <= "01000000"; -- 0x2a3
	when "01010100100" => qq <= "01001010"; -- 0x2a4
	when "01010100101" => qq <= "01001010"; -- 0x2a5
	when "01010100110" => qq <= "01001010"; -- 0x2a6
	when "01010100111" => qq <= "01001010"; -- 0x2a7
	when "01010101000" => qq <= "00101001"; -- 0x2a8
	when "01010101001" => qq <= "00001111"; -- 0x2a9
	when "01010101010" => qq <= "00000101"; -- 0x2aa
	when "01010101011" => qq <= "00101010"; -- 0x2ab
	when "01010101100" => qq <= "10000101"; -- 0x2ac
	when "01010101101" => qq <= "00101010"; -- 0x2ad
	when "01010101110" => qq <= "10100000"; -- 0x2ae
	when "01010101111" => qq <= "00000000"; -- 0x2af
	when "01010110000" => qq <= "10110001"; -- 0x2b0
	when "01010110001" => qq <= "00101000"; -- 0x2b1
	when "01010110010" => qq <= "11000101"; -- 0x2b2
	when "01010110011" => qq <= "00101010"; -- 0x2b3
	when "01010110100" => qq <= "11110000"; -- 0x2b4
	when "01010110101" => qq <= "00001000"; -- 0x2b5
	when "01010110110" => qq <= "11001000"; -- 0x2b6
	when "01010110111" => qq <= "11000000"; -- 0x2b7
	when "01010111000" => qq <= "00000100"; -- 0x2b8
	when "01010111001" => qq <= "11010000"; -- 0x2b9
	when "01010111010" => qq <= "11110101"; -- 0x2ba
	when "01010111011" => qq <= "01001100"; -- 0x2bb
	when "01010111100" => qq <= "00001010"; -- 0x2bc
	when "01010111101" => qq <= "00110011"; -- 0x2bd
	when "01010111110" => qq <= "10101101"; -- 0x2be
	when "01010111111" => qq <= "00101010"; -- 0x2bf
	when "01011000000" => qq <= "00000100"; -- 0x2c0
	when "01011000001" => qq <= "00011000"; -- 0x2c1
	when "01011000010" => qq <= "01101001"; -- 0x2c2
	when "01011000011" => qq <= "00000010"; -- 0x2c3
	when "01011000100" => qq <= "11001001"; -- 0x2c4
	when "01011000101" => qq <= "10111010"; -- 0x2c5
	when "01011000110" => qq <= "11010000"; -- 0x2c6
	when "01011000111" => qq <= "00011010"; -- 0x2c7
	when "01011001000" => qq <= "10101101"; -- 0x2c8
	when "01011001001" => qq <= "00101001"; -- 0x2c9
	when "01011001010" => qq <= "00000100"; -- 0x2ca
	when "01011001011" => qq <= "00011000"; -- 0x2cb
	when "01011001100" => qq <= "01101001"; -- 0x2cc
	when "01011001101" => qq <= "00000001"; -- 0x2cd
	when "01011001110" => qq <= "11001001"; -- 0x2ce
	when "01011001111" => qq <= "10111010"; -- 0x2cf
	when "01011010000" => qq <= "11010000"; -- 0x2d0
	when "01011010001" => qq <= "00001011"; -- 0x2d1
	when "01011010010" => qq <= "10101101"; -- 0x2d2
	when "01011010011" => qq <= "00101000"; -- 0x2d3
	when "01011010100" => qq <= "00000100"; -- 0x2d4
	when "01011010101" => qq <= "00011000"; -- 0x2d5
	when "01011010110" => qq <= "01101001"; -- 0x2d6
	when "01011010111" => qq <= "00000001"; -- 0x2d7
	when "01011011000" => qq <= "10001101"; -- 0x2d8
	when "01011011001" => qq <= "00101000"; -- 0x2d9
	when "01011011010" => qq <= "00000100"; -- 0x2da
	when "01011011011" => qq <= "10101001"; -- 0x2db
	when "01011011100" => qq <= "10110000"; -- 0x2dc
	when "01011011101" => qq <= "10001101"; -- 0x2dd
	when "01011011110" => qq <= "00101001"; -- 0x2de
	when "01011011111" => qq <= "00000100"; -- 0x2df
	when "01011100000" => qq <= "10101001"; -- 0x2e0
	when "01011100001" => qq <= "10110000"; -- 0x2e1
	when "01011100010" => qq <= "10001101"; -- 0x2e2
	when "01011100011" => qq <= "00101010"; -- 0x2e3
	when "01011100100" => qq <= "00000100"; -- 0x2e4
	when "01011100101" => qq <= "11001001"; -- 0x2e5
	when "01011100110" => qq <= "10110000"; -- 0x2e6
	when "01011100111" => qq <= "11010000"; -- 0x2e7
	when "01011101000" => qq <= "00100001"; -- 0x2e8
	when "01011101001" => qq <= "00101100"; -- 0x2e9
	when "01011101010" => qq <= "00110000"; -- 0x2ea
	when "01011101011" => qq <= "00001000"; -- 0x2eb
	when "01011101100" => qq <= "01110000"; -- 0x2ec
	when "01011101101" => qq <= "00001001"; -- 0x2ed
	when "01011101110" => qq <= "10100101"; -- 0x2ee
	when "01011101111" => qq <= "00110111"; -- 0x2ef
	when "01011110000" => qq <= "11010000"; -- 0x2f0
	when "01011110001" => qq <= "00000101"; -- 0x2f1
	when "01011110010" => qq <= "11100110"; -- 0x2f2
	when "01011110011" => qq <= "00110111"; -- 0x2f3
	when "01011110100" => qq <= "01001100"; -- 0x2f4
	when "01011110101" => qq <= "00001010"; -- 0x2f5
	when "01011110110" => qq <= "00110011"; -- 0x2f6
	when "01011110111" => qq <= "10101001"; -- 0x2f7
	when "01011111000" => qq <= "00000000"; -- 0x2f8
	when "01011111001" => qq <= "10000101"; -- 0x2f9
	when "01011111010" => qq <= "00110111"; -- 0x2fa
	when "01011111011" => qq <= "11100110"; -- 0x2fb
	when "01011111100" => qq <= "00110101"; -- 0x2fc
	when "01011111101" => qq <= "10100101"; -- 0x2fd
	when "01011111110" => qq <= "00110101"; -- 0x2fe
	when "01011111111" => qq <= "11001001"; -- 0x2ff
	when "01100000000" => qq <= "00001100"; -- 0x300
	when "01100000001" => qq <= "11010000"; -- 0x301
	when "01100000010" => qq <= "00000100"; -- 0x302
	when "01100000011" => qq <= "10101001"; -- 0x303
	when "01100000100" => qq <= "00000110"; -- 0x304
	when "01100000101" => qq <= "10000101"; -- 0x305
	when "01100000110" => qq <= "00110101"; -- 0x306
	when "01100000111" => qq <= "00100000"; -- 0x307
	when "01100001000" => qq <= "11001101"; -- 0x308
	when "01100001001" => qq <= "00111000"; -- 0x309
	when "01100001010" => qq <= "10100101"; -- 0x30a
	when "01100001011" => qq <= "00110001"; -- 0x30b
	when "01100001100" => qq <= "11110000"; -- 0x30c
	when "01100001101" => qq <= "00010101"; -- 0x30d
	when "01100001110" => qq <= "10100101"; -- 0x30e
	when "01100001111" => qq <= "00110000"; -- 0x30f
	when "01100010000" => qq <= "00101001"; -- 0x310
	when "01100010001" => qq <= "00100000"; -- 0x311
	when "01100010010" => qq <= "11110000"; -- 0x312
	when "01100010011" => qq <= "00001000"; -- 0x313
	when "01100010100" => qq <= "10100010"; -- 0x314
	when "01100010101" => qq <= "00000010"; -- 0x315
	when "01100010110" => qq <= "00100000"; -- 0x316
	when "01100010111" => qq <= "10110111"; -- 0x317
	when "01100011000" => qq <= "00111000"; -- 0x318
	when "01100011001" => qq <= "01001100"; -- 0x319
	when "01100011010" => qq <= "00100011"; -- 0x31a
	when "01100011011" => qq <= "00110011"; -- 0x31b
	when "01100011100" => qq <= "10100010"; -- 0x31c
	when "01100011101" => qq <= "00000010"; -- 0x31d
	when "01100011110" => qq <= "10101001"; -- 0x31e
	when "01100011111" => qq <= "00000000"; -- 0x31f
	when "01100100000" => qq <= "00100000"; -- 0x320
	when "01100100001" => qq <= "10001010"; -- 0x321
	when "01100100010" => qq <= "00111000"; -- 0x322
	when "01100100011" => qq <= "10101101"; -- 0x323
	when "01100100100" => qq <= "00101000"; -- 0x324
	when "01100100101" => qq <= "00000100"; -- 0x325
	when "01100100110" => qq <= "00101001"; -- 0x326
	when "01100100111" => qq <= "00111111"; -- 0x327
	when "01100101000" => qq <= "11000101"; -- 0x328
	when "01100101001" => qq <= "00111010"; -- 0x329
	when "01100101010" => qq <= "00110000"; -- 0x32a
	when "01100101011" => qq <= "00010011"; -- 0x32b
	when "01100101100" => qq <= "10101101"; -- 0x32c
	when "01100101101" => qq <= "00101001"; -- 0x32d
	when "01100101110" => qq <= "00000100"; -- 0x32e
	when "01100101111" => qq <= "00101001"; -- 0x32f
	when "01100110000" => qq <= "00111111"; -- 0x330
	when "01100110001" => qq <= "11000101"; -- 0x331
	when "01100110010" => qq <= "00111011"; -- 0x332
	when "01100110011" => qq <= "00110000"; -- 0x333
	when "01100110100" => qq <= "00001010"; -- 0x334
	when "01100110101" => qq <= "10100101"; -- 0x335
	when "01100110110" => qq <= "00110001"; -- 0x336
	when "01100110111" => qq <= "11010000"; -- 0x337
	when "01100111000" => qq <= "00000110"; -- 0x338
	when "01100111001" => qq <= "10100101"; -- 0x339
	when "01100111010" => qq <= "00110100"; -- 0x33a
	when "01100111011" => qq <= "11010000"; -- 0x33b
	when "01100111100" => qq <= "00000010"; -- 0x33c
	when "01100111101" => qq <= "11100110"; -- 0x33d
	when "01100111110" => qq <= "00110100"; -- 0x33e
	when "01100111111" => qq <= "11000110"; -- 0x33f
	when "01101000000" => qq <= "00111100"; -- 0x340
	when "01101000001" => qq <= "11010000"; -- 0x341
	when "01101000010" => qq <= "00110101"; -- 0x342
	when "01101000011" => qq <= "10100101"; -- 0x343
	when "01101000100" => qq <= "01010000"; -- 0x344
	when "01101000101" => qq <= "11010000"; -- 0x345
	when "01101000110" => qq <= "00010100"; -- 0x346
	when "01101000111" => qq <= "11100110"; -- 0x347
	when "01101001000" => qq <= "01010000"; -- 0x348
	when "01101001001" => qq <= "10101001"; -- 0x349
	when "01101001010" => qq <= "00100000"; -- 0x34a
	when "01101001011" => qq <= "10001101"; -- 0x34b
	when "01101001100" => qq <= "00111010"; -- 0x34c
	when "01101001101" => qq <= "00000100"; -- 0x34d
	when "01101001110" => qq <= "10101001"; -- 0x34e
	when "01101001111" => qq <= "10111001"; -- 0x34f
	when "01101010000" => qq <= "10001101"; -- 0x350
	when "01101010001" => qq <= "00111011"; -- 0x351
	when "01101010010" => qq <= "00000100"; -- 0x352
	when "01101010011" => qq <= "10101001"; -- 0x353
	when "01101010100" => qq <= "10111010"; -- 0x354
	when "01101010101" => qq <= "10001101"; -- 0x355
	when "01101010110" => qq <= "00111100"; -- 0x356
	when "01101010111" => qq <= "00000100"; -- 0x357
	when "01101011000" => qq <= "01001100"; -- 0x358
	when "01101011001" => qq <= "01110001"; -- 0x359
	when "01101011010" => qq <= "00110011"; -- 0x35a
	when "01101011011" => qq <= "10101101"; -- 0x35b
	when "01101011100" => qq <= "00111100"; -- 0x35c
	when "01101011101" => qq <= "00000100"; -- 0x35d
	when "01101011110" => qq <= "11001001"; -- 0x35e
	when "01101011111" => qq <= "10110000"; -- 0x35f
	when "01101100000" => qq <= "11010000"; -- 0x360
	when "01101100001" => qq <= "00001111"; -- 0x361
	when "01101100010" => qq <= "10101101"; -- 0x362
	when "01101100011" => qq <= "00111011"; -- 0x363
	when "01101100100" => qq <= "00000100"; -- 0x364
	when "01101100101" => qq <= "11001001"; -- 0x365
	when "01101100110" => qq <= "10110000"; -- 0x366
	when "01101100111" => qq <= "11110000"; -- 0x367
	when "01101101000" => qq <= "00010010"; -- 0x368
	when "01101101001" => qq <= "11001110"; -- 0x369
	when "01101101010" => qq <= "00111011"; -- 0x36a
	when "01101101011" => qq <= "00000100"; -- 0x36b
	when "01101101100" => qq <= "10101001"; -- 0x36c
	when "01101101101" => qq <= "10111010"; -- 0x36d
	when "01101101110" => qq <= "10001101"; -- 0x36e
	when "01101101111" => qq <= "00111100"; -- 0x36f
	when "01101110000" => qq <= "00000100"; -- 0x370
	when "01101110001" => qq <= "11001110"; -- 0x371
	when "01101110010" => qq <= "00111100"; -- 0x372
	when "01101110011" => qq <= "00000100"; -- 0x373
	when "01101110100" => qq <= "10100101"; -- 0x374
	when "01101110101" => qq <= "00111111"; -- 0x375
	when "01101110110" => qq <= "10000101"; -- 0x376
	when "01101110111" => qq <= "00111100"; -- 0x377
	when "01101111000" => qq <= "01001100"; -- 0x378
	when "01101111001" => qq <= "01101010"; -- 0x379
	when "01101111010" => qq <= "00110100"; -- 0x37a
	when "01101111011" => qq <= "10100101"; -- 0x37b
	when "01101111100" => qq <= "00110100"; -- 0x37c
	when "01101111101" => qq <= "11110000"; -- 0x37d
	when "01101111110" => qq <= "00011001"; -- 0x37e
	when "01101111111" => qq <= "10101001"; -- 0x37f
	when "01110000000" => qq <= "00000000"; -- 0x380
	when "01110000001" => qq <= "10000101"; -- 0x381
	when "01110000010" => qq <= "00110100"; -- 0x382
	when "01110000011" => qq <= "11100110"; -- 0x383
	when "01110000100" => qq <= "00110001"; -- 0x384
	when "01110000101" => qq <= "10101001"; -- 0x385
	when "01110000110" => qq <= "10110011"; -- 0x386
	when "01110000111" => qq <= "10001101"; -- 0x387
	when "01110001000" => qq <= "00111011"; -- 0x388
	when "01110001001" => qq <= "00000100"; -- 0x389
	when "01110001010" => qq <= "10101001"; -- 0x38a
	when "01110001011" => qq <= "00000000"; -- 0x38b
	when "01110001100" => qq <= "10100010"; -- 0x38c
	when "01110001101" => qq <= "00000010"; -- 0x38d
	when "01110001110" => qq <= "00100000"; -- 0x38e
	when "01110001111" => qq <= "10001010"; -- 0x38f
	when "01110010000" => qq <= "00111000"; -- 0x390
	when "01110010001" => qq <= "10100101"; -- 0x391
	when "01110010010" => qq <= "00111111"; -- 0x392
	when "01110010011" => qq <= "10000101"; -- 0x393
	when "01110010100" => qq <= "00111100"; -- 0x394
	when "01110010101" => qq <= "01001100"; -- 0x395
	when "01110010110" => qq <= "01101010"; -- 0x396
	when "01110010111" => qq <= "00110100"; -- 0x397
	when "01110011000" => qq <= "10001101"; -- 0x398
	when "01110011001" => qq <= "00000001"; -- 0x399
	when "01110011010" => qq <= "00001100"; -- 0x39a
	when "01110011011" => qq <= "10001101"; -- 0x39b
	when "01110011100" => qq <= "00010000"; -- 0x39c
	when "01110011101" => qq <= "00001100"; -- 0x39d
	when "01110011110" => qq <= "10101001"; -- 0x39e
	when "01110011111" => qq <= "00000000"; -- 0x39f
	when "01110100000" => qq <= "10000101"; -- 0x3a0
	when "01110100001" => qq <= "00010110"; -- 0x3a1
	when "01110100010" => qq <= "10000101"; -- 0x3a2
	when "01110100011" => qq <= "00010100"; -- 0x3a3
	when "01110100100" => qq <= "10100010"; -- 0x3a4
	when "01110100101" => qq <= "00000010"; -- 0x3a5
	when "01110100110" => qq <= "00100000"; -- 0x3a6
	when "01110100111" => qq <= "10110111"; -- 0x3a7
	when "01110101000" => qq <= "00111000"; -- 0x3a8
	when "01110101001" => qq <= "10100010"; -- 0x3a9
	when "01110101010" => qq <= "00001100"; -- 0x3aa
	when "01110101011" => qq <= "00100000"; -- 0x3ab
	when "01110101100" => qq <= "10110111"; -- 0x3ac
	when "01110101101" => qq <= "00111000"; -- 0x3ad
	when "01110101110" => qq <= "10101001"; -- 0x3ae
	when "01110101111" => qq <= "00000000"; -- 0x3af
	when "01110110000" => qq <= "10100010"; -- 0x3b0
	when "01110110001" => qq <= "00001100"; -- 0x3b1
	when "01110110010" => qq <= "00100000"; -- 0x3b2
	when "01110110011" => qq <= "10001010"; -- 0x3b3
	when "01110110100" => qq <= "00111000"; -- 0x3b4
	when "01110110101" => qq <= "10101001"; -- 0x3b5
	when "01110110110" => qq <= "00000000"; -- 0x3b6
	when "01110110111" => qq <= "10100010"; -- 0x3b7
	when "01110111000" => qq <= "00010110"; -- 0x3b8
	when "01110111001" => qq <= "00100000"; -- 0x3b9
	when "01110111010" => qq <= "10001010"; -- 0x3ba
	when "01110111011" => qq <= "00111000"; -- 0x3bb
	when "01110111100" => qq <= "10101101"; -- 0x3bc
	when "01110111101" => qq <= "00101000"; -- 0x3bd
	when "01110111110" => qq <= "00000100"; -- 0x3be
	when "01110111111" => qq <= "00101001"; -- 0x3bf
	when "01111000000" => qq <= "00001111"; -- 0x3c0
	when "01111000001" => qq <= "00001010"; -- 0x3c1
	when "01111000010" => qq <= "00001010"; -- 0x3c2
	when "01111000011" => qq <= "00001010"; -- 0x3c3
	when "01111000100" => qq <= "00001010"; -- 0x3c4
	when "01111000101" => qq <= "10000101"; -- 0x3c5
	when "01111000110" => qq <= "00100010"; -- 0x3c6
	when "01111000111" => qq <= "10101101"; -- 0x3c7
	when "01111001000" => qq <= "00101001"; -- 0x3c8
	when "01111001001" => qq <= "00000100"; -- 0x3c9
	when "01111001010" => qq <= "00101001"; -- 0x3ca
	when "01111001011" => qq <= "00001111"; -- 0x3cb
	when "01111001100" => qq <= "00000101"; -- 0x3cc
	when "01111001101" => qq <= "00100010"; -- 0x3cd
	when "01111001110" => qq <= "10000101"; -- 0x3ce
	when "01111001111" => qq <= "00100010"; -- 0x3cf
	when "01111010000" => qq <= "10100101"; -- 0x3d0
	when "01111010001" => qq <= "00100010"; -- 0x3d1
	when "01111010010" => qq <= "11000101"; -- 0x3d2
	when "01111010011" => qq <= "01010100"; -- 0x3d3
	when "01111010100" => qq <= "00110000"; -- 0x3d4
	when "01111010101" => qq <= "00000100"; -- 0x3d5
	when "01111010110" => qq <= "10100010"; -- 0x3d6
	when "01111010111" => qq <= "00011000"; -- 0x3d7
	when "01111011000" => qq <= "00010000"; -- 0x3d8
	when "01111011001" => qq <= "00001010"; -- 0x3d9
	when "01111011010" => qq <= "11000101"; -- 0x3da
	when "01111011011" => qq <= "01010101"; -- 0x3db
	when "01111011100" => qq <= "00110000"; -- 0x3dc
	when "01111011101" => qq <= "00000100"; -- 0x3dd
	when "01111011110" => qq <= "10100010"; -- 0x3de
	when "01111011111" => qq <= "00011010"; -- 0x3df
	when "01111100000" => qq <= "00010000"; -- 0x3e0
	when "01111100001" => qq <= "00000010"; -- 0x3e1
	when "01111100010" => qq <= "10100010"; -- 0x3e2
	when "01111100011" => qq <= "00011100"; -- 0x3e3
	when "01111100100" => qq <= "10101001"; -- 0x3e4
	when "01111100101" => qq <= "00000001"; -- 0x3e5
	when "01111100110" => qq <= "00100000"; -- 0x3e6
	when "01111100111" => qq <= "10001010"; -- 0x3e7
	when "01111101000" => qq <= "00111000"; -- 0x3e8
	when "01111101001" => qq <= "10100101"; -- 0x3e9
	when "01111101010" => qq <= "00100000"; -- 0x3ea
	when "01111101011" => qq <= "11010000"; -- 0x3eb
	when "01111101100" => qq <= "00000011"; -- 0x3ec
	when "01111101101" => qq <= "10001101"; -- 0x3ed
	when "01111101110" => qq <= "00110000"; -- 0x3ee
	when "01111101111" => qq <= "00001100"; -- 0x3ef
	when "01111110000" => qq <= "00100000"; -- 0x3f0
	when "01111110001" => qq <= "11101110"; -- 0x3f1
	when "01111110010" => qq <= "00111001"; -- 0x3f2
	when "01111110011" => qq <= "10101001"; -- 0x3f3
	when "01111110100" => qq <= "00001000"; -- 0x3f4
	when "01111110101" => qq <= "10100010"; -- 0x3f5
	when "01111110110" => qq <= "01111111"; -- 0x3f6
	when "01111110111" => qq <= "10100000"; -- 0x3f7
	when "01111111000" => qq <= "01111111"; -- 0x3f8
	when "01111111001" => qq <= "10000101"; -- 0x3f9
	when "01111111010" => qq <= "00100110"; -- 0x3fa
	when "01111111011" => qq <= "10000110"; -- 0x3fb
	when "01111111100" => qq <= "00101000"; -- 0x3fc
	when "01111111101" => qq <= "10000100"; -- 0x3fd
	when "01111111110" => qq <= "00101010"; -- 0x3fe
	when "01111111111" => qq <= "00100000"; -- 0x3ff
	when "10000000000" => qq <= "11111111"; -- 0x400
	when "10000000001" => qq <= "00110111"; -- 0x401
	when "10000000010" => qq <= "10100101"; -- 0x402
	when "10000000011" => qq <= "00110110"; -- 0x403
	when "10000000100" => qq <= "11010000"; -- 0x404
	when "10000000101" => qq <= "01001111"; -- 0x405
	when "10000000110" => qq <= "10100101"; -- 0x406
	when "10000000111" => qq <= "00100000"; -- 0x407
	when "10000001000" => qq <= "11110000"; -- 0x408
	when "10000001001" => qq <= "00001000"; -- 0x409
	when "10000001010" => qq <= "10001101"; -- 0x40a
	when "10000001011" => qq <= "00110001"; -- 0x40b
	when "10000001100" => qq <= "00001100"; -- 0x40c
	when "10000001101" => qq <= "00101100"; -- 0x40d
	when "10000001110" => qq <= "00101101"; -- 0x40e
	when "10000001111" => qq <= "00001000"; -- 0x40f
	when "10000010000" => qq <= "00010000"; -- 0x410
	when "10000010001" => qq <= "01000011"; -- 0x411
	when "10000010010" => qq <= "10100101"; -- 0x412
	when "10000010011" => qq <= "00100110"; -- 0x413
	when "10000010100" => qq <= "10100110"; -- 0x414
	when "10000010101" => qq <= "00101000"; -- 0x415
	when "10000010110" => qq <= "10100100"; -- 0x416
	when "10000010111" => qq <= "00101010"; -- 0x417
	when "10000011000" => qq <= "10001000"; -- 0x418
	when "10000011001" => qq <= "11010000"; -- 0x419
	when "10000011010" => qq <= "11011110"; -- 0x41a
	when "10000011011" => qq <= "10000101"; -- 0x41b
	when "10000011100" => qq <= "00101010"; -- 0x41c
	when "10000011101" => qq <= "10000110"; -- 0x41d
	when "10000011110" => qq <= "00101011"; -- 0x41e
	when "10000011111" => qq <= "11100110"; -- 0x41f
	when "10000100000" => qq <= "00110000"; -- 0x420
	when "10000100001" => qq <= "10100101"; -- 0x421
	when "10000100010" => qq <= "00110000"; -- 0x422
	when "10000100011" => qq <= "00101001"; -- 0x423
	when "10000100100" => qq <= "00100000"; -- 0x424
	when "10000100101" => qq <= "11110000"; -- 0x425
	when "10000100110" => qq <= "00001000"; -- 0x426
	when "10000100111" => qq <= "10100010"; -- 0x427
	when "10000101000" => qq <= "00010110"; -- 0x428
	when "10000101001" => qq <= "00100000"; -- 0x429
	when "10000101010" => qq <= "10110111"; -- 0x42a
	when "10000101011" => qq <= "00111000"; -- 0x42b
	when "10000101100" => qq <= "01001100"; -- 0x42c
	when "10000101101" => qq <= "00110110"; -- 0x42d
	when "10000101110" => qq <= "00110100"; -- 0x42e
	when "10000101111" => qq <= "10101001"; -- 0x42f
	when "10000110000" => qq <= "00000001"; -- 0x430
	when "10000110001" => qq <= "10100010"; -- 0x431
	when "10000110010" => qq <= "00010110"; -- 0x432
	when "10000110011" => qq <= "00100000"; -- 0x433
	when "10000110100" => qq <= "10001010"; -- 0x434
	when "10000110101" => qq <= "00111000"; -- 0x435
	when "10000110110" => qq <= "10100101"; -- 0x436
	when "10000110111" => qq <= "00101010"; -- 0x437
	when "10000111000" => qq <= "10100110"; -- 0x438
	when "10000111001" => qq <= "00101011"; -- 0x439
	when "10000111010" => qq <= "10001101"; -- 0x43a
	when "10000111011" => qq <= "10000000"; -- 0x43b
	when "10000111100" => qq <= "00001100"; -- 0x43c
	when "10000111101" => qq <= "10100000"; -- 0x43d
	when "10000111110" => qq <= "01111111"; -- 0x43e
	when "10000111111" => qq <= "11001010"; -- 0x43f
	when "10001000000" => qq <= "11010000"; -- 0x440
	when "10001000001" => qq <= "10110111"; -- 0x441
	when "10001000010" => qq <= "10100000"; -- 0x442
	when "10001000011" => qq <= "01111111"; -- 0x443
	when "10001000100" => qq <= "10100010"; -- 0x444
	when "10001000101" => qq <= "01111111"; -- 0x445
	when "10001000110" => qq <= "11001001"; -- 0x446
	when "10001000111" => qq <= "00001001"; -- 0x447
	when "10001001000" => qq <= "10010000"; -- 0x448
	when "10001001001" => qq <= "00000010"; -- 0x449
	when "10001001010" => qq <= "10101001"; -- 0x44a
	when "10001001011" => qq <= "00000101"; -- 0x44b
	when "10001001100" => qq <= "00111000"; -- 0x44c
	when "10001001101" => qq <= "11101001"; -- 0x44d
	when "10001001110" => qq <= "00000001"; -- 0x44e
	when "10001001111" => qq <= "00010000"; -- 0x44f
	when "10001010000" => qq <= "10101000"; -- 0x450
	when "10001010001" => qq <= "10101001"; -- 0x451
	when "10001010010" => qq <= "00000001"; -- 0x452
	when "10001010011" => qq <= "10000101"; -- 0x453
	when "10001010100" => qq <= "00101010"; -- 0x454
	when "10001010101" => qq <= "10100010"; -- 0x455
	when "10001010110" => qq <= "00010110"; -- 0x456
	when "10001010111" => qq <= "00100000"; -- 0x457
	when "10001011000" => qq <= "10110111"; -- 0x458
	when "10001011001" => qq <= "00111000"; -- 0x459
	when "10001011010" => qq <= "10100010"; -- 0x45a
	when "10001011011" => qq <= "00001100"; -- 0x45b
	when "10001011100" => qq <= "00100000"; -- 0x45c
	when "10001011101" => qq <= "10110111"; -- 0x45d
	when "10001011110" => qq <= "00111000"; -- 0x45e
	when "10001011111" => qq <= "10100101"; -- 0x45f
	when "10001100000" => qq <= "00100000"; -- 0x460
	when "10001100001" => qq <= "11010000"; -- 0x461
	when "10001100010" => qq <= "00000100"; -- 0x462
	when "10001100011" => qq <= "10001101"; -- 0x463
	when "10001100100" => qq <= "00110000"; -- 0x464
	when "10001100101" => qq <= "00001100"; -- 0x465
	when "10001100110" => qq <= "01100000"; -- 0x466
	when "10001100111" => qq <= "01001100"; -- 0x467
	when "10001101000" => qq <= "11111000"; -- 0x468
	when "10001101001" => qq <= "00110000"; -- 0x469
	when "10001101010" => qq <= "00100000"; -- 0x46a
	when "10001101011" => qq <= "11011000"; -- 0x46b
	when "10001101100" => qq <= "00110111"; -- 0x46c
	when "10001101101" => qq <= "00101100"; -- 0x46d
	when "10001101110" => qq <= "01000000"; -- 0x46e
	when "10001101111" => qq <= "00001000"; -- 0x46f
	when "10001110000" => qq <= "00010000"; -- 0x470
	when "10001110001" => qq <= "00000010"; -- 0x471
	when "10001110010" => qq <= "01110000"; -- 0x472
	when "10001110011" => qq <= "00000011"; -- 0x473
	when "10001110100" => qq <= "00100000"; -- 0x474
	when "10001110101" => qq <= "11111111"; -- 0x475
	when "10001110110" => qq <= "00110111"; -- 0x476
	when "10001110111" => qq <= "00101100"; -- 0x477
	when "10001111000" => qq <= "00000000"; -- 0x478
	when "10001111001" => qq <= "00001100"; -- 0x479
	when "10001111010" => qq <= "01010000"; -- 0x47a
	when "10001111011" => qq <= "11110001"; -- 0x47b
	when "10001111100" => qq <= "00100000"; -- 0x47c
	when "10001111101" => qq <= "00011011"; -- 0x47d
	when "10001111110" => qq <= "00110111"; -- 0x47e
	when "10001111111" => qq <= "10001101"; -- 0x47f
	when "10010000000" => qq <= "10000000"; -- 0x480
	when "10010000001" => qq <= "00001100"; -- 0x481
	when "10010000010" => qq <= "01001100"; -- 0x482
	when "10010000011" => qq <= "01011111"; -- 0x483
	when "10010000100" => qq <= "00110001"; -- 0x484
	when "10010000101" => qq <= "00100000"; -- 0x485
	when "10010000110" => qq <= "11001001"; -- 0x486
	when "10010000111" => qq <= "00110100"; -- 0x487
	when "10010001000" => qq <= "10110101"; -- 0x488
	when "10010001001" => qq <= "00000000"; -- 0x489
	when "10010001010" => qq <= "01001010"; -- 0x48a
	when "10010001011" => qq <= "01001010"; -- 0x48b
	when "10010001100" => qq <= "01001010"; -- 0x48c
	when "10010001101" => qq <= "01001010"; -- 0x48d
	when "10010001110" => qq <= "01001010"; -- 0x48e
	when "10010001111" => qq <= "00011000"; -- 0x48f
	when "10010010000" => qq <= "01101001"; -- 0x490
	when "10010010001" => qq <= "00000001"; -- 0x491
	when "10010010010" => qq <= "10000101"; -- 0x492
	when "10010010011" => qq <= "00100010"; -- 0x493
	when "10010010100" => qq <= "10100000"; -- 0x494
	when "10010010101" => qq <= "00000011"; -- 0x495
	when "10010010110" => qq <= "10110101"; -- 0x496
	when "10010010111" => qq <= "00000100"; -- 0x497
	when "10010011000" => qq <= "00111000"; -- 0x498
	when "10010011001" => qq <= "11110101"; -- 0x499
	when "10010011010" => qq <= "00101100"; -- 0x49a
	when "10010011011" => qq <= "00101001"; -- 0x49b
	when "10010011100" => qq <= "11111000"; -- 0x49c
	when "10010011101" => qq <= "11110000"; -- 0x49d
	when "10010011110" => qq <= "00010111"; -- 0x49e
	when "10010011111" => qq <= "00110000"; -- 0x49f
	when "10010100000" => qq <= "00000010"; -- 0x4a0
	when "10010100001" => qq <= "10100000"; -- 0x4a1
	when "10010100010" => qq <= "11111101"; -- 0x4a2
	when "10010100011" => qq <= "10011000"; -- 0x4a3
	when "10010100100" => qq <= "00011000"; -- 0x4a4
	when "10010100101" => qq <= "01110101"; -- 0x4a5
	when "10010100110" => qq <= "00000100"; -- 0x4a6
	when "10010100111" => qq <= "10010101"; -- 0x4a7
	when "10010101000" => qq <= "00000100"; -- 0x4a8
	when "10010101001" => qq <= "10000110"; -- 0x4a9
	when "10010101010" => qq <= "00100110"; -- 0x4aa
	when "10010101011" => qq <= "00000110"; -- 0x4ab
	when "10010101100" => qq <= "00100110"; -- 0x4ac
	when "10010101101" => qq <= "10100100"; -- 0x4ad
	when "10010101110" => qq <= "00100110"; -- 0x4ae
	when "10010101111" => qq <= "10011001"; -- 0x4af
	when "10010110000" => qq <= "00011001"; -- 0x4b0
	when "10010110001" => qq <= "00000000"; -- 0x4b1
	when "10010110010" => qq <= "10101001"; -- 0x4b2
	when "10010110011" => qq <= "11111111"; -- 0x4b3
	when "10010110100" => qq <= "10000101"; -- 0x4b4
	when "10010110101" => qq <= "00100010"; -- 0x4b5
	when "10010110110" => qq <= "10110101"; -- 0x4b6
	when "10010110111" => qq <= "00000000"; -- 0x4b7
	when "10010111000" => qq <= "00011000"; -- 0x4b8
	when "10010111001" => qq <= "01100101"; -- 0x4b9
	when "10010111010" => qq <= "00100010"; -- 0x4ba
	when "10010111011" => qq <= "11011101"; -- 0x4bb
	when "10010111100" => qq <= "10101001"; -- 0x4bc
	when "10010111101" => qq <= "00111100"; -- 0x4bd
	when "10010111110" => qq <= "10010000"; -- 0x4be
	when "10010111111" => qq <= "00000011"; -- 0x4bf
	when "10011000000" => qq <= "10111101"; -- 0x4c0
	when "10011000001" => qq <= "10101001"; -- 0x4c1
	when "10011000010" => qq <= "00111100"; -- 0x4c2
	when "10011000011" => qq <= "10010101"; -- 0x4c3
	when "10011000100" => qq <= "00000000"; -- 0x4c4
	when "10011000101" => qq <= "00100000"; -- 0x4c5
	when "10011000110" => qq <= "00010000"; -- 0x4c6
	when "10011000111" => qq <= "00110101"; -- 0x4c7
	when "10011001000" => qq <= "01100000"; -- 0x4c8
	when "10011001001" => qq <= "10101001"; -- 0x4c9
	when "10011001010" => qq <= "00000000"; -- 0x4ca
	when "10011001011" => qq <= "10000101"; -- 0x4cb
	when "10011001100" => qq <= "00100010"; -- 0x4cc
	when "10011001101" => qq <= "10101001"; -- 0x4cd
	when "10011001110" => qq <= "00000100"; -- 0x4ce
	when "10011001111" => qq <= "10000101"; -- 0x4cf
	when "10011010000" => qq <= "00100011"; -- 0x4d0
	when "10011010001" => qq <= "10110101"; -- 0x4d1
	when "10011010010" => qq <= "01000000"; -- 0x4d2
	when "10011010011" => qq <= "00011000"; -- 0x4d3
	when "10011010100" => qq <= "01101001"; -- 0x4d4
	when "10011010101" => qq <= "00000100"; -- 0x4d5
	when "10011010110" => qq <= "01001010"; -- 0x4d6
	when "10011010111" => qq <= "01001010"; -- 0x4d7
	when "10011011000" => qq <= "01001010"; -- 0x4d8
	when "10011011001" => qq <= "01001001"; -- 0x4d9
	when "10011011010" => qq <= "00011111"; -- 0x4da
	when "10011011011" => qq <= "00011000"; -- 0x4db
	when "10011011100" => qq <= "01100101"; -- 0x4dc
	when "10011011101" => qq <= "00100010"; -- 0x4dd
	when "10011011110" => qq <= "10000101"; -- 0x4de
	when "10011011111" => qq <= "00100010"; -- 0x4df
	when "10011100000" => qq <= "10101001"; -- 0x4e0
	when "10011100001" => qq <= "00000000"; -- 0x4e1
	when "10011100010" => qq <= "10000101"; -- 0x4e2
	when "10011100011" => qq <= "00100100"; -- 0x4e3
	when "10011100100" => qq <= "01100101"; -- 0x4e4
	when "10011100101" => qq <= "00100011"; -- 0x4e5
	when "10011100110" => qq <= "10000101"; -- 0x4e6
	when "10011100111" => qq <= "00100011"; -- 0x4e7
	when "10011101000" => qq <= "10110101"; -- 0x4e8
	when "10011101001" => qq <= "01000100"; -- 0x4e9
	when "10011101010" => qq <= "00011000"; -- 0x4ea
	when "10011101011" => qq <= "01101001"; -- 0x4eb
	when "10011101100" => qq <= "00000100"; -- 0x4ec
	when "10011101101" => qq <= "00001001"; -- 0x4ed
	when "10011101110" => qq <= "00000111"; -- 0x4ee
	when "10011101111" => qq <= "01001001"; -- 0x4ef
	when "10011110000" => qq <= "11111111"; -- 0x4f0
	when "10011110001" => qq <= "00001010"; -- 0x4f1
	when "10011110010" => qq <= "00100110"; -- 0x4f2
	when "10011110011" => qq <= "00100100"; -- 0x4f3
	when "10011110100" => qq <= "00001010"; -- 0x4f4
	when "10011110101" => qq <= "00100110"; -- 0x4f5
	when "10011110110" => qq <= "00100100"; -- 0x4f6
	when "10011110111" => qq <= "00011000"; -- 0x4f7
	when "10011111000" => qq <= "01100101"; -- 0x4f8
	when "10011111001" => qq <= "00100010"; -- 0x4f9
	when "10011111010" => qq <= "10000101"; -- 0x4fa
	when "10011111011" => qq <= "00100010"; -- 0x4fb
	when "10011111100" => qq <= "10100101"; -- 0x4fc
	when "10011111101" => qq <= "00100100"; -- 0x4fd
	when "10011111110" => qq <= "01100101"; -- 0x4fe
	when "10011111111" => qq <= "00100011"; -- 0x4ff
	when "10100000000" => qq <= "10000101"; -- 0x500
	when "10100000001" => qq <= "00100011"; -- 0x501
	when "10100000010" => qq <= "10100000"; -- 0x502
	when "10100000011" => qq <= "00000000"; -- 0x503
	when "10100000100" => qq <= "10110001"; -- 0x504
	when "10100000101" => qq <= "00100010"; -- 0x505
	when "10100000110" => qq <= "00010000"; -- 0x506
	when "10100000111" => qq <= "00000111"; -- 0x507
	when "10100001000" => qq <= "00001010"; -- 0x508
	when "10100001001" => qq <= "00001010"; -- 0x509
	when "10100001010" => qq <= "00001010"; -- 0x50a
	when "10100001011" => qq <= "00001010"; -- 0x50b
	when "10100001100" => qq <= "00001010"; -- 0x50c
	when "10100001101" => qq <= "10010101"; -- 0x50d
	when "10100001110" => qq <= "00101100"; -- 0x50e
	when "10100001111" => qq <= "01100000"; -- 0x50f
	when "10100010000" => qq <= "10000110"; -- 0x510
	when "10100010001" => qq <= "00100010"; -- 0x511
	when "10100010010" => qq <= "10101001"; -- 0x512
	when "10100010011" => qq <= "00000000"; -- 0x513
	when "10100010100" => qq <= "10000101"; -- 0x514
	when "10100010101" => qq <= "01010010"; -- 0x515
	when "10100010110" => qq <= "10110101"; -- 0x516
	when "10100010111" => qq <= "00000000"; -- 0x517
	when "10100011000" => qq <= "11110000"; -- 0x518
	when "10100011001" => qq <= "01110010"; -- 0x519
	when "10100011010" => qq <= "01001010"; -- 0x51a
	when "10100011011" => qq <= "01001010"; -- 0x51b
	when "10100011100" => qq <= "01001010"; -- 0x51c
	when "10100011101" => qq <= "10000101"; -- 0x51d
	when "10100011110" => qq <= "00100100"; -- 0x51e
	when "10100011111" => qq <= "10110101"; -- 0x51f
	when "10100100000" => qq <= "00000100"; -- 0x520
	when "10100100001" => qq <= "01001010"; -- 0x521
	when "10100100010" => qq <= "01001010"; -- 0x522
	when "10100100011" => qq <= "01001010"; -- 0x523
	when "10100100100" => qq <= "10101010"; -- 0x524
	when "10100100101" => qq <= "10000110"; -- 0x525
	when "10100100110" => qq <= "00100110"; -- 0x526
	when "10100100111" => qq <= "10111101"; -- 0x527
	when "10100101000" => qq <= "00000110"; -- 0x528
	when "10100101001" => qq <= "00101111"; -- 0x529
	when "10100101010" => qq <= "11110000"; -- 0x52a
	when "10100101011" => qq <= "00101101"; -- 0x52b
	when "10100101100" => qq <= "00001010"; -- 0x52c
	when "10100101101" => qq <= "10101010"; -- 0x52d
	when "10100101110" => qq <= "00100000"; -- 0x52e
	when "10100101111" => qq <= "10100111"; -- 0x52f
	when "10100110000" => qq <= "00110101"; -- 0x530
	when "10100110001" => qq <= "10100110"; -- 0x531
	when "10100110010" => qq <= "00100010"; -- 0x532
	when "10100110011" => qq <= "10100101"; -- 0x533
	when "10100110100" => qq <= "00101000"; -- 0x534
	when "10100110101" => qq <= "00011000"; -- 0x535
	when "10100110110" => qq <= "01110101"; -- 0x536
	when "10100110111" => qq <= "00001000"; -- 0x537
	when "10100111000" => qq <= "10010101"; -- 0x538
	when "10100111001" => qq <= "00001000"; -- 0x539
	when "10100111010" => qq <= "10100101"; -- 0x53a
	when "10100111011" => qq <= "00101001"; -- 0x53b
	when "10100111100" => qq <= "01110101"; -- 0x53c
	when "10100111101" => qq <= "01000000"; -- 0x53d
	when "10100111110" => qq <= "00010000"; -- 0x53e
	when "10100111111" => qq <= "00010111"; -- 0x53f
	when "10101000000" => qq <= "11001001"; -- 0x540
	when "10101000001" => qq <= "11111100"; -- 0x541
	when "10101000010" => qq <= "00110000"; -- 0x542
	when "10101000011" => qq <= "00001000"; -- 0x543
	when "10101000100" => qq <= "10101001"; -- 0x544
	when "10101000101" => qq <= "00000001"; -- 0x545
	when "10101000110" => qq <= "10000101"; -- 0x546
	when "10101000111" => qq <= "01010010"; -- 0x547
	when "10101001000" => qq <= "10101001"; -- 0x548
	when "10101001001" => qq <= "00000000"; -- 0x549
	when "10101001010" => qq <= "11110000"; -- 0x54a
	when "10101001011" => qq <= "00001011"; -- 0x54b
	when "10101001100" => qq <= "11001001"; -- 0x54c
	when "10101001101" => qq <= "11110111"; -- 0x54d
	when "10101001110" => qq <= "00110000"; -- 0x54e
	when "10101001111" => qq <= "00000111"; -- 0x54f
	when "10101010000" => qq <= "10101001"; -- 0x550
	when "10101010001" => qq <= "00000001"; -- 0x551
	when "10101010010" => qq <= "10001101"; -- 0x552
	when "10101010011" => qq <= "01010010"; -- 0x553
	when "10101010100" => qq <= "00000000"; -- 0x554
	when "10101010101" => qq <= "10101001"; -- 0x555
	when "10101010110" => qq <= "11110111"; -- 0x556
	when "10101010111" => qq <= "10010101"; -- 0x557
	when "10101011000" => qq <= "01000000"; -- 0x558
	when "10101011001" => qq <= "10100110"; -- 0x559
	when "10101011010" => qq <= "00100110"; -- 0x55a
	when "10101011011" => qq <= "10111101"; -- 0x55b
	when "10101011100" => qq <= "00100110"; -- 0x55c
	when "10101011101" => qq <= "00101111"; -- 0x55d
	when "10101011110" => qq <= "11110000"; -- 0x55e
	when "10101011111" => qq <= "00101100"; -- 0x55f
	when "10101100000" => qq <= "00001010"; -- 0x560
	when "10101100001" => qq <= "10101010"; -- 0x561
	when "10101100010" => qq <= "00100000"; -- 0x562
	when "10101100011" => qq <= "10100111"; -- 0x563
	when "10101100100" => qq <= "00110101"; -- 0x564
	when "10101100101" => qq <= "10100110"; -- 0x565
	when "10101100110" => qq <= "00100010"; -- 0x566
	when "10101100111" => qq <= "10100101"; -- 0x567
	when "10101101000" => qq <= "00101000"; -- 0x568
	when "10101101001" => qq <= "00011000"; -- 0x569
	when "10101101010" => qq <= "01110101"; -- 0x56a
	when "10101101011" => qq <= "00001100"; -- 0x56b
	when "10101101100" => qq <= "10010101"; -- 0x56c
	when "10101101101" => qq <= "00001100"; -- 0x56d
	when "10101101110" => qq <= "10100101"; -- 0x56e
	when "10101101111" => qq <= "00101001"; -- 0x56f
	when "10101110000" => qq <= "01110101"; -- 0x570
	when "10101110001" => qq <= "01000100"; -- 0x571
	when "10101110010" => qq <= "00010000"; -- 0x572
	when "10101110011" => qq <= "00001100"; -- 0x573
	when "10101110100" => qq <= "11001001"; -- 0x574
	when "10101110101" => qq <= "11101000"; -- 0x575
	when "10101110110" => qq <= "00110000"; -- 0x576
	when "10101110111" => qq <= "00010010"; -- 0x577
	when "10101111000" => qq <= "10101001"; -- 0x578
	when "10101111001" => qq <= "00000001"; -- 0x579
	when "10101111010" => qq <= "10000101"; -- 0x57a
	when "10101111011" => qq <= "01010010"; -- 0x57b
	when "10101111100" => qq <= "10101001"; -- 0x57c
	when "10101111101" => qq <= "11101000"; -- 0x57d
	when "10101111110" => qq <= "00110000"; -- 0x57e
	when "10101111111" => qq <= "00001010"; -- 0x57f
	when "10110000000" => qq <= "11001001"; -- 0x580
	when "10110000001" => qq <= "00100000"; -- 0x581
	when "10110000010" => qq <= "00010000"; -- 0x582
	when "10110000011" => qq <= "00000110"; -- 0x583
	when "10110000100" => qq <= "10101001"; -- 0x584
	when "10110000101" => qq <= "00000001"; -- 0x585
	when "10110000110" => qq <= "10000101"; -- 0x586
	when "10110000111" => qq <= "01010010"; -- 0x587
	when "10110001000" => qq <= "10101001"; -- 0x588
	when "10110001001" => qq <= "00100000"; -- 0x589
	when "10110001010" => qq <= "10010101"; -- 0x58a
	when "10110001011" => qq <= "01000100"; -- 0x58b
	when "10110001100" => qq <= "10100110"; -- 0x58c
	when "10110001101" => qq <= "00100010"; -- 0x58d
	when "10110001110" => qq <= "11100000"; -- 0x58e
	when "10110001111" => qq <= "00000000"; -- 0x58f
	when "10110010000" => qq <= "11110000"; -- 0x590
	when "10110010001" => qq <= "00010100"; -- 0x591
	when "10110010010" => qq <= "10100101"; -- 0x592
	when "10110010011" => qq <= "01010010"; -- 0x593
	when "10110010100" => qq <= "11110000"; -- 0x594
	when "10110010101" => qq <= "00010000"; -- 0x595
	when "10110010110" => qq <= "10101001"; -- 0x596
	when "10110010111" => qq <= "00100000"; -- 0x597
	when "10110011000" => qq <= "10010101"; -- 0x598
	when "10110011001" => qq <= "01000000"; -- 0x599
	when "10110011010" => qq <= "10101001"; -- 0x59a
	when "10110011011" => qq <= "01010000"; -- 0x59b
	when "10110011100" => qq <= "10010101"; -- 0x59c
	when "10110011101" => qq <= "01000100"; -- 0x59d
	when "10110011110" => qq <= "10101001"; -- 0x59e
	when "10110011111" => qq <= "11000000"; -- 0x59f
	when "10110100000" => qq <= "10010101"; -- 0x5a0
	when "10110100001" => qq <= "00000100"; -- 0x5a1
	when "10110100010" => qq <= "10101001"; -- 0x5a2
	when "10110100011" => qq <= "00000001"; -- 0x5a3
	when "10110100100" => qq <= "10010101"; -- 0x5a4
	when "10110100101" => qq <= "00000000"; -- 0x5a5
	when "10110100110" => qq <= "01100000"; -- 0x5a6
	when "10110100111" => qq <= "10000110"; -- 0x5a7
	when "10110101000" => qq <= "00100101"; -- 0x5a8
	when "10110101001" => qq <= "10001010"; -- 0x5a9
	when "10110101010" => qq <= "00010000"; -- 0x5aa
	when "10110101011" => qq <= "00000110"; -- 0x5ab
	when "10110101100" => qq <= "01001001"; -- 0x5ac
	when "10110101101" => qq <= "11111111"; -- 0x5ad
	when "10110101110" => qq <= "00011000"; -- 0x5ae
	when "10110101111" => qq <= "01101001"; -- 0x5af
	when "10110110000" => qq <= "00000001"; -- 0x5b0
	when "10110110001" => qq <= "10101010"; -- 0x5b1
	when "10110110010" => qq <= "10101001"; -- 0x5b2
	when "10110110011" => qq <= "00000000"; -- 0x5b3
	when "10110110100" => qq <= "10000101"; -- 0x5b4
	when "10110110101" => qq <= "00101000"; -- 0x5b5
	when "10110110110" => qq <= "10000101"; -- 0x5b6
	when "10110110111" => qq <= "00101001"; -- 0x5b7
	when "10110111000" => qq <= "10100101"; -- 0x5b8
	when "10110111001" => qq <= "00101000"; -- 0x5b9
	when "10110111010" => qq <= "00011000"; -- 0x5ba
	when "10110111011" => qq <= "01100101"; -- 0x5bb
	when "10110111100" => qq <= "00100100"; -- 0x5bc
	when "10110111101" => qq <= "10000101"; -- 0x5bd
	when "10110111110" => qq <= "00101000"; -- 0x5be
	when "10110111111" => qq <= "10101001"; -- 0x5bf
	when "10111000000" => qq <= "00000000"; -- 0x5c0
	when "10111000001" => qq <= "01100101"; -- 0x5c1
	when "10111000010" => qq <= "00101001"; -- 0x5c2
	when "10111000011" => qq <= "10000101"; -- 0x5c3
	when "10111000100" => qq <= "00101001"; -- 0x5c4
	when "10111000101" => qq <= "11001010"; -- 0x5c5
	when "10111000110" => qq <= "11010000"; -- 0x5c6
	when "10111000111" => qq <= "11110000"; -- 0x5c7
	when "10111001000" => qq <= "10100101"; -- 0x5c8
	when "10111001001" => qq <= "00100101"; -- 0x5c9
	when "10111001010" => qq <= "00010000"; -- 0x5ca
	when "10111001011" => qq <= "00001101"; -- 0x5cb
	when "10111001100" => qq <= "10101001"; -- 0x5cc
	when "10111001101" => qq <= "00000000"; -- 0x5cd
	when "10111001110" => qq <= "00111000"; -- 0x5ce
	when "10111001111" => qq <= "11100101"; -- 0x5cf
	when "10111010000" => qq <= "00101000"; -- 0x5d0
	when "10111010001" => qq <= "10000101"; -- 0x5d1
	when "10111010010" => qq <= "00101000"; -- 0x5d2
	when "10111010011" => qq <= "10101001"; -- 0x5d3
	when "10111010100" => qq <= "00000000"; -- 0x5d4
	when "10111010101" => qq <= "11100101"; -- 0x5d5
	when "10111010110" => qq <= "00101001"; -- 0x5d6
	when "10111010111" => qq <= "10000101"; -- 0x5d7
	when "10111011000" => qq <= "00101001"; -- 0x5d8
	when "10111011001" => qq <= "01100000"; -- 0x5d9
	when "10111011010" => qq <= "10100010"; -- 0x5da
	when "10111011011" => qq <= "00000000"; -- 0x5db
	when "10111011100" => qq <= "10101001"; -- 0x5dc
	when "10111011101" => qq <= "00100000"; -- 0x5dd
	when "10111011110" => qq <= "10100000"; -- 0x5de
	when "10111011111" => qq <= "00000000"; -- 0x5df
	when "10111100000" => qq <= "10010101"; -- 0x5e0
	when "10111100001" => qq <= "01000000"; -- 0x5e1
	when "10111100010" => qq <= "10010100"; -- 0x5e2
	when "10111100011" => qq <= "00001000"; -- 0x5e3
	when "10111100100" => qq <= "10010100"; -- 0x5e4
	when "10111100101" => qq <= "00001100"; -- 0x5e5
	when "10111100110" => qq <= "11101000"; -- 0x5e6
	when "10111100111" => qq <= "11100000"; -- 0x5e7
	when "10111101000" => qq <= "00000100"; -- 0x5e8
	when "10111101001" => qq <= "11010000"; -- 0x5e9
	when "10111101010" => qq <= "11110101"; -- 0x5ea
	when "10111101011" => qq <= "10100010"; -- 0x5eb
	when "10111101100" => qq <= "00000000"; -- 0x5ec
	when "10111101101" => qq <= "10101001"; -- 0x5ed
	when "10111101110" => qq <= "00000001"; -- 0x5ee
	when "10111101111" => qq <= "10010101"; -- 0x5ef
	when "10111110000" => qq <= "00000000"; -- 0x5f0
	when "10111110001" => qq <= "11101000"; -- 0x5f1
	when "10111110010" => qq <= "11100000"; -- 0x5f2
	when "10111110011" => qq <= "00000100"; -- 0x5f3
	when "10111110100" => qq <= "11010000"; -- 0x5f4
	when "10111110101" => qq <= "11111001"; -- 0x5f5
	when "10111110110" => qq <= "10100010"; -- 0x5f6
	when "10111110111" => qq <= "00000000"; -- 0x5f7
	when "10111111000" => qq <= "10100000"; -- 0x5f8
	when "10111111001" => qq <= "00000000"; -- 0x5f9
	when "10111111010" => qq <= "10101001"; -- 0x5fa
	when "10111111011" => qq <= "11000000"; -- 0x5fb
	when "10111111100" => qq <= "10010101"; -- 0x5fc
	when "10111111101" => qq <= "00000100"; -- 0x5fd
	when "10111111110" => qq <= "10011001"; -- 0x5fe
	when "10111111111" => qq <= "00011001"; -- 0x5ff
	when "11000000000" => qq <= "00000000"; -- 0x600
	when "11000000001" => qq <= "11001000"; -- 0x601
	when "11000000010" => qq <= "11001000"; -- 0x602
	when "11000000011" => qq <= "11101000"; -- 0x603
	when "11000000100" => qq <= "11100000"; -- 0x604
	when "11000000101" => qq <= "00000100"; -- 0x605
	when "11000000110" => qq <= "11010000"; -- 0x606
	when "11000000111" => qq <= "11110100"; -- 0x607
	when "11000001000" => qq <= "10101001"; -- 0x608
	when "11000001001" => qq <= "01010000"; -- 0x609
	when "11000001010" => qq <= "10000101"; -- 0x60a
	when "11000001011" => qq <= "01000100"; -- 0x60b
	when "11000001100" => qq <= "10101001"; -- 0x60c
	when "11000001101" => qq <= "01000100"; -- 0x60d
	when "11000001110" => qq <= "10000101"; -- 0x60e
	when "11000001111" => qq <= "01000101"; -- 0x60f
	when "11000010000" => qq <= "10101001"; -- 0x610
	when "11000010001" => qq <= "00111000"; -- 0x611
	when "11000010010" => qq <= "10000101"; -- 0x612
	when "11000010011" => qq <= "01000110"; -- 0x613
	when "11000010100" => qq <= "10101001"; -- 0x614
	when "11000010101" => qq <= "00101100"; -- 0x615
	when "11000010110" => qq <= "10000101"; -- 0x616
	when "11000010111" => qq <= "01000111"; -- 0x617
	when "11000011000" => qq <= "10101101"; -- 0x618
	when "11000011001" => qq <= "00110011"; -- 0x619
	when "11000011010" => qq <= "00001000"; -- 0x61a
	when "11000011011" => qq <= "01001001"; -- 0x61b
	when "11000011100" => qq <= "11111111"; -- 0x61c
	when "11000011101" => qq <= "00011000"; -- 0x61d
	when "11000011110" => qq <= "00101010"; -- 0x61e
	when "11000011111" => qq <= "00101010"; -- 0x61f
	when "11000100000" => qq <= "00101010"; -- 0x620
	when "11000100001" => qq <= "00101001"; -- 0x621
	when "11000100010" => qq <= "00000011"; -- 0x622
	when "11000100011" => qq <= "10101000"; -- 0x623
	when "11000100100" => qq <= "10111001"; -- 0x624
	when "11000100101" => qq <= "10100101"; -- 0x625
	when "11000100110" => qq <= "00111100"; -- 0x626
	when "11000100111" => qq <= "10000101"; -- 0x627
	when "11000101000" => qq <= "00111100"; -- 0x628
	when "11000101001" => qq <= "10000101"; -- 0x629
	when "11000101010" => qq <= "00111111"; -- 0x62a
	when "11000101011" => qq <= "10101001"; -- 0x62b
	when "11000101100" => qq <= "00000100"; -- 0x62c
	when "11000101101" => qq <= "10000101"; -- 0x62d
	when "11000101110" => qq <= "01010100"; -- 0x62e
	when "11000101111" => qq <= "10101001"; -- 0x62f
	when "11000110000" => qq <= "00000010"; -- 0x630
	when "11000110001" => qq <= "10000101"; -- 0x631
	when "11000110010" => qq <= "01010101"; -- 0x632
	when "11000110011" => qq <= "10101001"; -- 0x633
	when "11000110100" => qq <= "00000011"; -- 0x634
	when "11000110101" => qq <= "10000101"; -- 0x635
	when "11000110110" => qq <= "01010110"; -- 0x636
	when "11000110111" => qq <= "10101101"; -- 0x637
	when "11000111000" => qq <= "00110011"; -- 0x638
	when "11000111001" => qq <= "00001000"; -- 0x639
	when "11000111010" => qq <= "01001001"; -- 0x63a
	when "11000111011" => qq <= "11111111"; -- 0x63b
	when "11000111100" => qq <= "00011000"; -- 0x63c
	when "11000111101" => qq <= "00101010"; -- 0x63d
	when "11000111110" => qq <= "00101010"; -- 0x63e
	when "11000111111" => qq <= "00101010"; -- 0x63f
	when "11001000000" => qq <= "00101001"; -- 0x640
	when "11001000001" => qq <= "00000011"; -- 0x641
	when "11001000010" => qq <= "00011000"; -- 0x642
	when "11001000011" => qq <= "01101001"; -- 0x643
	when "11001000100" => qq <= "00000010"; -- 0x644
	when "11001000101" => qq <= "10000101"; -- 0x645
	when "11001000110" => qq <= "00100010"; -- 0x646
	when "11001000111" => qq <= "10100010"; -- 0x647
	when "11001001000" => qq <= "00000000"; -- 0x648
	when "11001001001" => qq <= "10000110"; -- 0x649
	when "11001001010" => qq <= "00100100"; -- 0x64a
	when "11001001011" => qq <= "10000110"; -- 0x64b
	when "11001001100" => qq <= "00100110"; -- 0x64c
	when "11001001101" => qq <= "10000110"; -- 0x64d
	when "11001001110" => qq <= "00101000"; -- 0x64e
	when "11001001111" => qq <= "10100101"; -- 0x64f
	when "11001010000" => qq <= "00100100"; -- 0x650
	when "11001010001" => qq <= "11111000"; -- 0x651
	when "11001010010" => qq <= "00011000"; -- 0x652
	when "11001010011" => qq <= "01100101"; -- 0x653
	when "11001010100" => qq <= "01010100"; -- 0x654
	when "11001010101" => qq <= "10000101"; -- 0x655
	when "11001010110" => qq <= "00100100"; -- 0x656
	when "11001010111" => qq <= "10100101"; -- 0x657
	when "11001011000" => qq <= "00100110"; -- 0x658
	when "11001011001" => qq <= "00011000"; -- 0x659
	when "11001011010" => qq <= "01100101"; -- 0x65a
	when "11001011011" => qq <= "01010101"; -- 0x65b
	when "11001011100" => qq <= "10000101"; -- 0x65c
	when "11001011101" => qq <= "00100110"; -- 0x65d
	when "11001011110" => qq <= "10100101"; -- 0x65e
	when "11001011111" => qq <= "00101000"; -- 0x65f
	when "11001100000" => qq <= "00011000"; -- 0x660
	when "11001100001" => qq <= "01100101"; -- 0x661
	when "11001100010" => qq <= "01010110"; -- 0x662
	when "11001100011" => qq <= "10000101"; -- 0x663
	when "11001100100" => qq <= "00101000"; -- 0x664
	when "11001100101" => qq <= "11011000"; -- 0x665
	when "11001100110" => qq <= "11101000"; -- 0x666
	when "11001100111" => qq <= "11100100"; -- 0x667
	when "11001101000" => qq <= "00100010"; -- 0x668
	when "11001101001" => qq <= "11010000"; -- 0x669
	when "11001101010" => qq <= "11100100"; -- 0x66a
	when "11001101011" => qq <= "10100101"; -- 0x66b
	when "11001101100" => qq <= "00100100"; -- 0x66c
	when "11001101101" => qq <= "10000101"; -- 0x66d
	when "11001101110" => qq <= "01010100"; -- 0x66e
	when "11001101111" => qq <= "10100101"; -- 0x66f
	when "11001110000" => qq <= "00100110"; -- 0x670
	when "11001110001" => qq <= "10000101"; -- 0x671
	when "11001110010" => qq <= "01010101"; -- 0x672
	when "11001110011" => qq <= "10100101"; -- 0x673
	when "11001110100" => qq <= "00101000"; -- 0x674
	when "11001110101" => qq <= "10000101"; -- 0x675
	when "11001110110" => qq <= "01010110"; -- 0x676
	when "11001110111" => qq <= "10101101"; -- 0x677
	when "11001111000" => qq <= "00110010"; -- 0x678
	when "11001111001" => qq <= "00001000"; -- 0x679
	when "11001111010" => qq <= "00010000"; -- 0x67a
	when "11001111011" => qq <= "00001101"; -- 0x67b
	when "11001111100" => qq <= "10101001"; -- 0x67c
	when "11001111101" => qq <= "01000000"; -- 0x67d
	when "11001111110" => qq <= "10000101"; -- 0x67e
	when "11001111111" => qq <= "00111010"; -- 0x67f
	when "11010000000" => qq <= "10000101"; -- 0x680
	when "11010000001" => qq <= "00111011"; -- 0x681
	when "11010000010" => qq <= "10100101"; -- 0x682
	when "11010000011" => qq <= "01010110"; -- 0x683
	when "11010000100" => qq <= "10000101"; -- 0x684
	when "11010000101" => qq <= "01010100"; -- 0x685
	when "11010000110" => qq <= "01001100"; -- 0x686
	when "11010000111" => qq <= "10011101"; -- 0x687
	when "11010001000" => qq <= "00110110"; -- 0x688
	when "11010001001" => qq <= "10100101"; -- 0x689
	when "11010001010" => qq <= "01010110"; -- 0x68a
	when "11010001011" => qq <= "00101001"; -- 0x68b
	when "11010001100" => qq <= "11110000"; -- 0x68c
	when "11010001101" => qq <= "01001010"; -- 0x68d
	when "11010001110" => qq <= "01001010"; -- 0x68e
	when "11010001111" => qq <= "01001010"; -- 0x68f
	when "11010010000" => qq <= "01001010"; -- 0x690
	when "11010010001" => qq <= "00001001"; -- 0x691
	when "11010010010" => qq <= "00110000"; -- 0x692
	when "11010010011" => qq <= "10000101"; -- 0x693
	when "11010010100" => qq <= "00111010"; -- 0x694
	when "11010010101" => qq <= "10100101"; -- 0x695
	when "11010010110" => qq <= "01010110"; -- 0x696
	when "11010010111" => qq <= "00101001"; -- 0x697
	when "11010011000" => qq <= "00001111"; -- 0x698
	when "11010011001" => qq <= "00001001"; -- 0x699
	when "11010011010" => qq <= "00110000"; -- 0x69a
	when "11010011011" => qq <= "10000101"; -- 0x69b
	when "11010011100" => qq <= "00111011"; -- 0x69c
	when "11010011101" => qq <= "10101001"; -- 0x69d
	when "11010011110" => qq <= "00000000"; -- 0x69e
	when "11010011111" => qq <= "10000101"; -- 0x69f
	when "11010100000" => qq <= "00110111"; -- 0x6a0
	when "11010100001" => qq <= "10000101"; -- 0x6a1
	when "11010100010" => qq <= "00110000"; -- 0x6a2
	when "11010100011" => qq <= "10001101"; -- 0x6a3
	when "11010100100" => qq <= "00010000"; -- 0x6a4
	when "11010100101" => qq <= "00001100"; -- 0x6a5
	when "11010100110" => qq <= "10000101"; -- 0x6a6
	when "11010100111" => qq <= "00010100"; -- 0x6a7
	when "11010101000" => qq <= "10000101"; -- 0x6a8
	when "11010101001" => qq <= "00010101"; -- 0x6a9
	when "11010101010" => qq <= "10000101"; -- 0x6aa
	when "11010101011" => qq <= "00110011"; -- 0x6ab
	when "11010101100" => qq <= "10000101"; -- 0x6ac
	when "11010101101" => qq <= "00111101"; -- 0x6ad
	when "11010101110" => qq <= "10000101"; -- 0x6ae
	when "11010101111" => qq <= "00111110"; -- 0x6af
	when "11010110000" => qq <= "10000101"; -- 0x6b0
	when "11010110001" => qq <= "00111000"; -- 0x6b1
	when "11010110010" => qq <= "10000101"; -- 0x6b2
	when "11010110011" => qq <= "00110100"; -- 0x6b3
	when "11010110100" => qq <= "10000101"; -- 0x6b4
	when "11010110101" => qq <= "00110001"; -- 0x6b5
	when "11010110110" => qq <= "10000101"; -- 0x6b6
	when "11010110111" => qq <= "01010000"; -- 0x6b7
	when "11010111000" => qq <= "10001101"; -- 0x6b8
	when "11010111001" => qq <= "00010110"; -- 0x6b9
	when "11010111010" => qq <= "00000000"; -- 0x6ba
	when "11010111011" => qq <= "10001101"; -- 0x6bb
	when "11010111100" => qq <= "00000000"; -- 0x6bc
	when "11010111101" => qq <= "00001101"; -- 0x6bd
	when "11010111110" => qq <= "10001101"; -- 0x6be
	when "11010111111" => qq <= "00000000"; -- 0x6bf
	when "11011000000" => qq <= "00001110"; -- 0x6c0
	when "11011000001" => qq <= "10101101"; -- 0x6c1
	when "11011000010" => qq <= "00101010"; -- 0x6c2
	when "11011000011" => qq <= "00000100"; -- 0x6c3
	when "11011000100" => qq <= "10000101"; -- 0x6c4
	when "11011000101" => qq <= "00100110"; -- 0x6c5
	when "11011000110" => qq <= "10101101"; -- 0x6c6
	when "11011000111" => qq <= "00101001"; -- 0x6c7
	when "11011001000" => qq <= "00000100"; -- 0x6c8
	when "11011001001" => qq <= "10000101"; -- 0x6c9
	when "11011001010" => qq <= "00100111"; -- 0x6ca
	when "11011001011" => qq <= "10101101"; -- 0x6cb
	when "11011001100" => qq <= "00101000"; -- 0x6cc
	when "11011001101" => qq <= "00000100"; -- 0x6cd
	when "11011001110" => qq <= "10000101"; -- 0x6ce
	when "11011001111" => qq <= "00101011"; -- 0x6cf
	when "11011010000" => qq <= "10101001"; -- 0x6d0
	when "11011010001" => qq <= "00000001"; -- 0x6d1
	when "11011010010" => qq <= "10100010"; -- 0x6d2
	when "11011010011" => qq <= "00000100"; -- 0x6d3
	when "11011010100" => qq <= "00100000"; -- 0x6d4
	when "11011010101" => qq <= "10001010"; -- 0x6d5
	when "11011010110" => qq <= "00111000"; -- 0x6d6
	when "11011010111" => qq <= "10100101"; -- 0x6d7
	when "11011011000" => qq <= "00100110"; -- 0x6d8
	when "11011011001" => qq <= "10001101"; -- 0x6d9
	when "11011011010" => qq <= "00101010"; -- 0x6da
	when "11011011011" => qq <= "00000100"; -- 0x6db
	when "11011011100" => qq <= "10100101"; -- 0x6dc
	when "11011011101" => qq <= "00100111"; -- 0x6dd
	when "11011011110" => qq <= "10001101"; -- 0x6de
	when "11011011111" => qq <= "00101001"; -- 0x6df
	when "11011100000" => qq <= "00000100"; -- 0x6e0
	when "11011100001" => qq <= "10100101"; -- 0x6e1
	when "11011100010" => qq <= "00101011"; -- 0x6e2
	when "11011100011" => qq <= "10001101"; -- 0x6e3
	when "11011100100" => qq <= "00101000"; -- 0x6e4
	when "11011100101" => qq <= "00000100"; -- 0x6e5
	when "11011100110" => qq <= "10100101"; -- 0x6e6
	when "11011100111" => qq <= "00101010"; -- 0x6e7
	when "11011101000" => qq <= "11010000"; -- 0x6e8
	when "11011101001" => qq <= "00001011"; -- 0x6e9
	when "11011101010" => qq <= "10101001"; -- 0x6ea
	when "11011101011" => qq <= "10110000"; -- 0x6eb
	when "11011101100" => qq <= "10001101"; -- 0x6ec
	when "11011101101" => qq <= "00101010"; -- 0x6ed
	when "11011101110" => qq <= "00000100"; -- 0x6ee
	when "11011101111" => qq <= "10001101"; -- 0x6ef
	when "11011110000" => qq <= "00101001"; -- 0x6f0
	when "11011110001" => qq <= "00000100"; -- 0x6f1
	when "11011110010" => qq <= "10001101"; -- 0x6f2
	when "11011110011" => qq <= "00101000"; -- 0x6f3
	when "11011110100" => qq <= "00000100"; -- 0x6f4
	when "11011110101" => qq <= "10101001"; -- 0x6f5
	when "11011110110" => qq <= "10110000"; -- 0x6f6
	when "11011110111" => qq <= "10001101"; -- 0x6f7
	when "11011111000" => qq <= "00111011"; -- 0x6f8
	when "11011111001" => qq <= "00000100"; -- 0x6f9
	when "11011111010" => qq <= "10001101"; -- 0x6fa
	when "11011111011" => qq <= "00111100"; -- 0x6fb
	when "11011111100" => qq <= "00000100"; -- 0x6fc
	when "11011111101" => qq <= "10101001"; -- 0x6fd
	when "11011111110" => qq <= "10110001"; -- 0x6fe
	when "11011111111" => qq <= "10001101"; -- 0x6ff
	when "11100000000" => qq <= "00111010"; -- 0x700
	when "11100000001" => qq <= "00000100"; -- 0x701
	when "11100000010" => qq <= "01100000"; -- 0x702
	when "11100000011" => qq <= "10101001"; -- 0x703
	when "11100000100" => qq <= "00000000"; -- 0x704
	when "11100000101" => qq <= "10000101"; -- 0x705
	when "11100000110" => qq <= "00100000"; -- 0x706
	when "11100000111" => qq <= "10000101"; -- 0x707
	when "11100001000" => qq <= "00110110"; -- 0x708
	when "11100001001" => qq <= "10001101"; -- 0x709
	when "11100001010" => qq <= "00110000"; -- 0x70a
	when "11100001011" => qq <= "00001100"; -- 0x70b
	when "11100001100" => qq <= "10000101"; -- 0x70c
	when "11100001101" => qq <= "00101010"; -- 0x70d
	when "11100001110" => qq <= "10101001"; -- 0x70e
	when "11100001111" => qq <= "00110000"; -- 0x70f
	when "11100010000" => qq <= "10000101"; -- 0x710
	when "11100010001" => qq <= "01010111"; -- 0x711
	when "11100010010" => qq <= "10000101"; -- 0x712
	when "11100010011" => qq <= "01011000"; -- 0x713
	when "11100010100" => qq <= "10000101"; -- 0x714
	when "11100010101" => qq <= "01011001"; -- 0x715
	when "11100010110" => qq <= "10101001"; -- 0x716
	when "11100010111" => qq <= "00000110"; -- 0x717
	when "11100011000" => qq <= "10000101"; -- 0x718
	when "11100011001" => qq <= "01010001"; -- 0x719
	when "11100011010" => qq <= "01100000"; -- 0x71a
	when "11100011011" => qq <= "10101101"; -- 0x71b
	when "11100011100" => qq <= "00101010"; -- 0x71c
	when "11100011101" => qq <= "00000100"; -- 0x71d
	when "11100011110" => qq <= "00101001"; -- 0x71e
	when "11100011111" => qq <= "00111111"; -- 0x71f
	when "11100100000" => qq <= "00100000"; -- 0x720
	when "11100100001" => qq <= "01110001"; -- 0x721
	when "11100100010" => qq <= "00110111"; -- 0x722
	when "11100100011" => qq <= "10100101"; -- 0x723
	when "11100100100" => qq <= "00100010"; -- 0x724
	when "11100100101" => qq <= "11110000"; -- 0x725
	when "11100100110" => qq <= "00000101"; -- 0x726
	when "11100100111" => qq <= "10101001"; -- 0x727
	when "11100101000" => qq <= "10110000"; -- 0x728
	when "11100101001" => qq <= "10001101"; -- 0x729
	when "11100101010" => qq <= "00101010"; -- 0x72a
	when "11100101011" => qq <= "00000100"; -- 0x72b
	when "11100101100" => qq <= "10101101"; -- 0x72c
	when "11100101101" => qq <= "00101001"; -- 0x72d
	when "11100101110" => qq <= "00000100"; -- 0x72e
	when "11100101111" => qq <= "00101001"; -- 0x72f
	when "11100110000" => qq <= "00111111"; -- 0x730
	when "11100110001" => qq <= "00100000"; -- 0x731
	when "11100110010" => qq <= "01110001"; -- 0x732
	when "11100110011" => qq <= "00110111"; -- 0x733
	when "11100110100" => qq <= "10100101"; -- 0x734
	when "11100110101" => qq <= "00100010"; -- 0x735
	when "11100110110" => qq <= "11110000"; -- 0x736
	when "11100110111" => qq <= "00000101"; -- 0x737
	when "11100111000" => qq <= "10101001"; -- 0x738
	when "11100111001" => qq <= "10110000"; -- 0x739
	when "11100111010" => qq <= "10001101"; -- 0x73a
	when "11100111011" => qq <= "00101001"; -- 0x73b
	when "11100111100" => qq <= "00000100"; -- 0x73c
	when "11100111101" => qq <= "10101101"; -- 0x73d
	when "11100111110" => qq <= "00101000"; -- 0x73e
	when "11100111111" => qq <= "00000100"; -- 0x73f
	when "11101000000" => qq <= "00101001"; -- 0x740
	when "11101000001" => qq <= "00111111"; -- 0x741
	when "11101000010" => qq <= "00100000"; -- 0x742
	when "11101000011" => qq <= "01110001"; -- 0x743
	when "11101000100" => qq <= "00110111"; -- 0x744
	when "11101000101" => qq <= "10100101"; -- 0x745
	when "11101000110" => qq <= "00100010"; -- 0x746
	when "11101000111" => qq <= "11110000"; -- 0x747
	when "11101001000" => qq <= "00000101"; -- 0x748
	when "11101001001" => qq <= "10101001"; -- 0x749
	when "11101001010" => qq <= "10110000"; -- 0x74a
	when "11101001011" => qq <= "10001101"; -- 0x74b
	when "11101001100" => qq <= "00101000"; -- 0x74c
	when "11101001101" => qq <= "00000100"; -- 0x74d
	when "11101001110" => qq <= "10101101"; -- 0x74e
	when "11101001111" => qq <= "00111011"; -- 0x74f
	when "11101010000" => qq <= "00000100"; -- 0x750
	when "11101010001" => qq <= "00101001"; -- 0x751
	when "11101010010" => qq <= "00111111"; -- 0x752
	when "11101010011" => qq <= "00100000"; -- 0x753
	when "11101010100" => qq <= "01110001"; -- 0x754
	when "11101010101" => qq <= "00110111"; -- 0x755
	when "11101010110" => qq <= "10100101"; -- 0x756
	when "11101010111" => qq <= "00100010"; -- 0x757
	when "11101011000" => qq <= "11110000"; -- 0x758
	when "11101011001" => qq <= "00000101"; -- 0x759
	when "11101011010" => qq <= "10101001"; -- 0x75a
	when "11101011011" => qq <= "10111001"; -- 0x75b
	when "11101011100" => qq <= "10001101"; -- 0x75c
	when "11101011101" => qq <= "00111011"; -- 0x75d
	when "11101011110" => qq <= "00000100"; -- 0x75e
	when "11101011111" => qq <= "10101101"; -- 0x75f
	when "11101100000" => qq <= "00111100"; -- 0x760
	when "11101100001" => qq <= "00000100"; -- 0x761
	when "11101100010" => qq <= "00101001"; -- 0x762
	when "11101100011" => qq <= "00111111"; -- 0x763
	when "11101100100" => qq <= "00100000"; -- 0x764
	when "11101100101" => qq <= "01110001"; -- 0x765
	when "11101100110" => qq <= "00110111"; -- 0x766
	when "11101100111" => qq <= "10100101"; -- 0x767
	when "11101101000" => qq <= "00100010"; -- 0x768
	when "11101101001" => qq <= "11110000"; -- 0x769
	when "11101101010" => qq <= "00000101"; -- 0x76a
	when "11101101011" => qq <= "10101001"; -- 0x76b
	when "11101101100" => qq <= "10111001"; -- 0x76c
	when "11101101101" => qq <= "10001101"; -- 0x76d
	when "11101101110" => qq <= "00111100"; -- 0x76e
	when "11101101111" => qq <= "00000100"; -- 0x76f
	when "11101110000" => qq <= "01100000"; -- 0x770
	when "11101110001" => qq <= "11001001"; -- 0x771
	when "11101110010" => qq <= "00110000"; -- 0x772
	when "11101110011" => qq <= "10010000"; -- 0x773
	when "11101110100" => qq <= "00001000"; -- 0x774
	when "11101110101" => qq <= "11001001"; -- 0x775
	when "11101110110" => qq <= "00111010"; -- 0x776
	when "11101110111" => qq <= "10110000"; -- 0x777
	when "11101111000" => qq <= "00000100"; -- 0x778
	when "11101111001" => qq <= "10101001"; -- 0x779
	when "11101111010" => qq <= "00000000"; -- 0x77a
	when "11101111011" => qq <= "11110000"; -- 0x77b
	when "11101111100" => qq <= "00000010"; -- 0x77c
	when "11101111101" => qq <= "10101001"; -- 0x77d
	when "11101111110" => qq <= "00000001"; -- 0x77e
	when "11101111111" => qq <= "10000101"; -- 0x77f
	when "11110000000" => qq <= "00100010"; -- 0x780
	when "11110000001" => qq <= "01100000"; -- 0x781
	when "11110000010" => qq <= "10000110"; -- 0x782
	when "11110000011" => qq <= "00100110"; -- 0x783
	when "11110000100" => qq <= "10101001"; -- 0x784
	when "11110000101" => qq <= "00000000"; -- 0x785
	when "11110000110" => qq <= "10000101"; -- 0x786
	when "11110000111" => qq <= "00110010"; -- 0x787
	when "11110001000" => qq <= "00101100"; -- 0x788
	when "11110001001" => qq <= "00101000"; -- 0x789
	when "11110001010" => qq <= "00001000"; -- 0x78a
	when "11110001011" => qq <= "00010000"; -- 0x78b
	when "11110001100" => qq <= "00010000"; -- 0x78c
	when "11110001101" => qq <= "11100110"; -- 0x78d
	when "11110001110" => qq <= "00110010"; -- 0x78e
	when "11110001111" => qq <= "00101100"; -- 0x78f
	when "11110010000" => qq <= "00101001"; -- 0x790
	when "11110010001" => qq <= "00001000"; -- 0x791
	when "11110010010" => qq <= "00010000"; -- 0x792
	when "11110010011" => qq <= "00001001"; -- 0x793
	when "11110010100" => qq <= "11100110"; -- 0x794
	when "11110010101" => qq <= "00110010"; -- 0x795
	when "11110010110" => qq <= "00101100"; -- 0x796
	when "11110010111" => qq <= "00101010"; -- 0x797
	when "11110011000" => qq <= "00001000"; -- 0x798
	when "11110011001" => qq <= "00010000"; -- 0x799
	when "11110011010" => qq <= "00000010"; -- 0x79a
	when "11110011011" => qq <= "11100110"; -- 0x79b
	when "11110011100" => qq <= "00110010"; -- 0x79c
	when "11110011101" => qq <= "10110101"; -- 0x79d
	when "11110011110" => qq <= "00000000"; -- 0x79e
	when "11110011111" => qq <= "00101001"; -- 0x79f
	when "11110100000" => qq <= "11111000"; -- 0x7a0
	when "11110100001" => qq <= "01001010"; -- 0x7a1
	when "11110100010" => qq <= "01001010"; -- 0x7a2
	when "11110100011" => qq <= "10101010"; -- 0x7a3
	when "11110100100" => qq <= "10101001"; -- 0x7a4
	when "11110100101" => qq <= "00000010"; -- 0x7a5
	when "11110100110" => qq <= "00100100"; -- 0x7a6
	when "11110100111" => qq <= "00110010"; -- 0x7a7
	when "11110101000" => qq <= "11110000"; -- 0x7a8
	when "11110101001" => qq <= "00000001"; -- 0x7a9
	when "11110101010" => qq <= "11101000"; -- 0x7aa
	when "11110101011" => qq <= "10111101"; -- 0x7ab
	when "11110101100" => qq <= "01000110"; -- 0x7ac
	when "11110101101" => qq <= "00101111"; -- 0x7ad
	when "11110101110" => qq <= "00101100"; -- 0x7ae
	when "11110101111" => qq <= "00101011"; -- 0x7af
	when "11110110000" => qq <= "00001000"; -- 0x7b0
	when "11110110001" => qq <= "00110000"; -- 0x7b1
	when "11110110010" => qq <= "00000011"; -- 0x7b2
	when "11110110011" => qq <= "10111101"; -- 0x7b3
	when "11110110100" => qq <= "10000110"; -- 0x7b4
	when "11110110101" => qq <= "00101111"; -- 0x7b5
	when "11110110110" => qq <= "00011000"; -- 0x7b6
	when "11110110111" => qq <= "01000110"; -- 0x7b7
	when "11110111000" => qq <= "00110010"; -- 0x7b8
	when "11110111001" => qq <= "10110000"; -- 0x7b9
	when "11110111010" => qq <= "00000110"; -- 0x7ba
	when "11110111011" => qq <= "00101001"; -- 0x7bb
	when "11110111100" => qq <= "11110000"; -- 0x7bc
	when "11110111101" => qq <= "01001010"; -- 0x7bd
	when "11110111110" => qq <= "01001010"; -- 0x7be
	when "11110111111" => qq <= "01001010"; -- 0x7bf
	when "11111000000" => qq <= "01001010"; -- 0x7c0
	when "11111000001" => qq <= "00101001"; -- 0x7c1
	when "11111000010" => qq <= "00001111"; -- 0x7c2
	when "11111000011" => qq <= "10000101"; -- 0x7c3
	when "11111000100" => qq <= "00100100"; -- 0x7c4
	when "11111000101" => qq <= "00100110"; -- 0x7c5
	when "11111000110" => qq <= "00110010"; -- 0x7c6
	when "11111000111" => qq <= "10101001"; -- 0x7c7
	when "11111001000" => qq <= "00001000"; -- 0x7c8
	when "11111001001" => qq <= "00100100"; -- 0x7c9
	when "11111001010" => qq <= "00100100"; -- 0x7ca
	when "11111001011" => qq <= "11110000"; -- 0x7cb
	when "11111001100" => qq <= "00000110"; -- 0x7cc
	when "11111001101" => qq <= "10100101"; -- 0x7cd
	when "11111001110" => qq <= "00100100"; -- 0x7ce
	when "11111001111" => qq <= "00001001"; -- 0x7cf
	when "11111010000" => qq <= "11110000"; -- 0x7d0
	when "11111010001" => qq <= "10000101"; -- 0x7d1
	when "11111010010" => qq <= "00100100"; -- 0x7d2
	when "11111010011" => qq <= "10100101"; -- 0x7d3
	when "11111010100" => qq <= "00100100"; -- 0x7d4
	when "11111010101" => qq <= "10100110"; -- 0x7d5
	when "11111010110" => qq <= "00100110"; -- 0x7d6
	when "11111010111" => qq <= "01100000"; -- 0x7d7
	when "11111011000" => qq <= "10100010"; -- 0x7d8
	when "11111011001" => qq <= "00000000"; -- 0x7d9
	when "11111011010" => qq <= "10100000"; -- 0x7da
	when "11111011011" => qq <= "00000000"; -- 0x7db
	when "11111011100" => qq <= "10100101"; -- 0x7dc
	when "11111011101" => qq <= "00110011"; -- 0x7dd
	when "11111011110" => qq <= "11010000"; -- 0x7de
	when "11111011111" => qq <= "00011110"; -- 0x7df
	when "11111100000" => qq <= "00101100"; -- 0x7e0
	when "11111100001" => qq <= "10000000"; -- 0x7e1
	when "11111100010" => qq <= "00001000"; -- 0x7e2
	when "11111100011" => qq <= "00110000"; -- 0x7e3
	when "11111100100" => qq <= "00011001"; -- 0x7e4
	when "11111100101" => qq <= "10101001"; -- 0x7e5
	when "11111100110" => qq <= "00000011"; -- 0x7e6
	when "11111100111" => qq <= "10000101"; -- 0x7e7
	when "11111101000" => qq <= "00100010"; -- 0x7e8
	when "11111101001" => qq <= "00101100"; -- 0x7e9
	when "11111101010" => qq <= "10000000"; -- 0x7ea
	when "11111101011" => qq <= "00001000"; -- 0x7eb
	when "11111101100" => qq <= "01110000"; -- 0x7ec
	when "11111101101" => qq <= "00000100"; -- 0x7ed
	when "11111101110" => qq <= "10101001"; -- 0x7ee
	when "11111101111" => qq <= "11111101"; -- 0x7ef
	when "11111110000" => qq <= "10000101"; -- 0x7f0
	when "11111110001" => qq <= "00100010"; -- 0x7f1
	when "11111110010" => qq <= "10111001"; -- 0x7f2
	when "11111110011" => qq <= "00011001"; -- 0x7f3
	when "11111110100" => qq <= "00000000"; -- 0x7f4
	when "11111110101" => qq <= "00011000"; -- 0x7f5
	when "11111110110" => qq <= "01100101"; -- 0x7f6
	when "11111110111" => qq <= "00100010"; -- 0x7f7
	when "11111111000" => qq <= "10011001"; -- 0x7f8
	when "11111111001" => qq <= "00011001"; -- 0x7f9
	when "11111111010" => qq <= "00000000"; -- 0x7fa
	when "11111111011" => qq <= "10001101"; -- 0x7fb
	when "11111111100" => qq <= "00000000"; -- 0x7fc
	when "11111111101" => qq <= "00001110"; -- 0x7fd
	when "11111111110" => qq <= "01100000"; -- 0x7fe
	when "11111111111" => qq <= "00100000"; -- 0x7ff
	when others => qq <= "00000000";
END CASE; 
END PROCESS; 
END SYN; 
