module prog_rom4(input clock,
	input [10:0] address,
	output [7:0] q
	);

	reg [7:0] qq;
always @(posedge clk )
		case (address)
	13'h000: qq = 8'h30; // 0x000
	13'h001: qq = 8'h38; // 0x001
	13'h002: qq = 8'ha9; // 0x002
	13'h003: qq = 8'h0a; // 0x003
	13'h004: qq = 8'h85; // 0x004
	13'h005: qq = 8'h51; // 0x005
	13'h006: qq = 8'h2c; // 0x006
	13'h007: qq = 8'h31; // 0x007
	13'h008: qq = 8'h08; // 0x008
	13'h009: qq = 8'h10; // 0x009
	13'h00a: qq = 8'h11; // 0x00a
	13'h00b: qq = 8'h70; // 0x00b
	13'h00c: qq = 8'h1e; // 0x00c
	13'h00d: qq = 8'ha9; // 0x00d
	13'h00e: qq = 8'h08; // 0x00e
	13'h00f: qq = 8'h85; // 0x00f
	13'h010: qq = 8'h51; // 0x010
	13'h011: qq = 8'ha5; // 0x011
	13'h012: qq = 8'h36; // 0x012
	13'h013: qq = 8'hc9; // 0x013
	13'h014: qq = 8'h02; // 0x014
	13'h015: qq = 8'hf0; // 0x015
	13'h016: qq = 8'h01; // 0x016
	13'h017: qq = 8'h60; // 0x017
	13'h018: qq = 8'hc6; // 0x018
	13'h019: qq = 8'h36; // 0x019
	13'h01a: qq = 8'h10; // 0x01a
	13'h01b: qq = 8'h0f; // 0x01b
	13'h01c: qq = 8'h70; // 0x01c
	13'h01d: qq = 8'h04; // 0x01d
	13'h01e: qq = 8'ha9; // 0x01e
	13'h01f: qq = 8'h06; // 0x01f
	13'h020: qq = 8'h85; // 0x020
	13'h021: qq = 8'h51; // 0x021
	13'h022: qq = 8'ha5; // 0x022
	13'h023: qq = 8'h36; // 0x023
	13'h024: qq = 8'hd0; // 0x024
	13'h025: qq = 8'h01; // 0x025
	13'h026: qq = 8'h60; // 0x026
	13'h027: qq = 8'h50; // 0x027
	13'h028: qq = 8'h02; // 0x028
	13'h029: qq = 8'he6; // 0x029
	13'h02a: qq = 8'h20; // 0x02a
	13'h02b: qq = 8'he6; // 0x02b
	13'h02c: qq = 8'h20; // 0x02c
	13'h02d: qq = 8'hc6; // 0x02d
	13'h02e: qq = 8'h36; // 0x02e
	13'h02f: qq = 8'h60; // 0x02f
	13'h030: qq = 8'ha9; // 0x030
	13'h031: qq = 8'h09; // 0x031
	13'h032: qq = 8'h85; // 0x032
	13'h033: qq = 8'h22; // 0x033
	13'h034: qq = 8'h85; // 0x034
	13'h035: qq = 8'h23; // 0x035
	13'h036: qq = 8'h85; // 0x036
	13'h037: qq = 8'h24; // 0x037
	13'h038: qq = 8'h85; // 0x038
	13'h039: qq = 8'h25; // 0x039
	13'h03a: qq = 8'h2c; // 0x03a
	13'h03b: qq = 8'h40; // 0x03b
	13'h03c: qq = 8'h08; // 0x03c
	13'h03d: qq = 8'h10; // 0x03d
	13'h03e: qq = 8'h0b; // 0x03e
	13'h03f: qq = 8'h50; // 0x03f
	13'h040: qq = 8'h09; // 0x040
	13'h041: qq = 8'ha5; // 0x041
	13'h042: qq = 8'h22; // 0x042
	13'h043: qq = 8'h25; // 0x043
	13'h044: qq = 8'h23; // 0x044
	13'h045: qq = 8'hc9; // 0x045
	13'h046: qq = 8'h09; // 0x046
	13'h047: qq = 8'hd0; // 0x047
	13'h048: qq = 8'h01; // 0x048
	13'h049: qq = 8'h60; // 0x049
	13'h04a: qq = 8'h8d; // 0x04a
	13'h04b: qq = 8'h80; // 0x04b
	13'h04c: qq = 8'h0c; // 0x04c
	13'h04d: qq = 8'ha2; // 0x04d
	13'h04e: qq = 8'h01; // 0x04e
	13'h04f: qq = 8'ha0; // 0x04f
	13'h050: qq = 8'hfa; // 0x050
	13'h051: qq = 8'h88; // 0x051
	13'h052: qq = 8'hd0; // 0x052
	13'h053: qq = 8'hfd; // 0x053
	13'h054: qq = 8'h8a; // 0x054
	13'h055: qq = 8'hd0; // 0x055
	13'h056: qq = 8'h07; // 0x056
	13'h057: qq = 8'h2c; // 0x057
	13'h058: qq = 8'h40; // 0x058
	13'h059: qq = 8'h08; // 0x059
	13'h05a: qq = 8'h50; // 0x05a
	13'h05b: qq = 8'h1f; // 0x05b
	13'h05c: qq = 8'h70; // 0x05c
	13'h05d: qq = 8'h05; // 0x05d
	13'h05e: qq = 8'h2c; // 0x05e
	13'h05f: qq = 8'h40; // 0x05f
	13'h060: qq = 8'h08; // 0x060
	13'h061: qq = 8'h10; // 0x061
	13'h062: qq = 8'h18; // 0x062
	13'h063: qq = 8'hb5; // 0x063
	13'h064: qq = 8'h22; // 0x064
	13'h065: qq = 8'hf0; // 0x065
	13'h066: qq = 8'h06; // 0x066
	13'h067: qq = 8'ha9; // 0x067
	13'h068: qq = 8'h09; // 0x068
	13'h069: qq = 8'h95; // 0x069
	13'h06a: qq = 8'h22; // 0x06a
	13'h06b: qq = 8'hd0; // 0x06b
	13'h06c: qq = 8'h18; // 0x06c
	13'h06d: qq = 8'hd6; // 0x06d
	13'h06e: qq = 8'h24; // 0x06e
	13'h06f: qq = 8'hd0; // 0x06f
	13'h070: qq = 8'h14; // 0x070
	13'h071: qq = 8'he6; // 0x071
	13'h072: qq = 8'h36; // 0x072
	13'h073: qq = 8'ha9; // 0x073
	13'h074: qq = 8'h09; // 0x074
	13'h075: qq = 8'h95; // 0x075
	13'h076: qq = 8'h22; // 0x076
	13'h077: qq = 8'h95; // 0x077
	13'h078: qq = 8'h24; // 0x078
	13'h079: qq = 8'hd0; // 0x079
	13'h07a: qq = 8'h0a; // 0x07a
	13'h07b: qq = 8'ha9; // 0x07b
	13'h07c: qq = 8'h09; // 0x07c
	13'h07d: qq = 8'h95; // 0x07d
	13'h07e: qq = 8'h24; // 0x07e
	13'h07f: qq = 8'hb5; // 0x07f
	13'h080: qq = 8'h22; // 0x080
	13'h081: qq = 8'hf0; // 0x081
	13'h082: qq = 8'h02; // 0x082
	13'h083: qq = 8'hd6; // 0x083
	13'h084: qq = 8'h22; // 0x084
	13'h085: qq = 8'hca; // 0x085
	13'h086: qq = 8'h10; // 0x086
	13'h087: qq = 8'hcc; // 0x087
	13'h088: qq = 8'h30; // 0x088
	13'h089: qq = 8'hb0; // 0x089
	13'h08a: qq = 8'ha0; // 0x08a
	13'h08b: qq = 8'h00; // 0x08b
	13'h08c: qq = 8'hc9; // 0x08c
	13'h08d: qq = 8'h00; // 0x08d
	13'h08e: qq = 8'hf0; // 0x08e
	13'h08f: qq = 8'h02; // 0x08f
	13'h090: qq = 8'ha0; // 0x090
	13'h091: qq = 8'h80; // 0x091
	13'h092: qq = 8'h84; // 0x092
	13'h093: qq = 8'h28; // 0x093
	13'h094: qq = 8'hbd; // 0x094
	13'h095: qq = 8'h4f; // 0x095
	13'h096: qq = 8'h3c; // 0x096
	13'h097: qq = 8'h85; // 0x097
	13'h098: qq = 8'h22; // 0x098
	13'h099: qq = 8'hbd; // 0x099
	13'h09a: qq = 8'h50; // 0x09a
	13'h09b: qq = 8'h3c; // 0x09b
	13'h09c: qq = 8'h85; // 0x09c
	13'h09d: qq = 8'h23; // 0x09d
	13'h09e: qq = 8'hbd; // 0x09e
	13'h09f: qq = 8'h71; // 0x09f
	13'h0a0: qq = 8'h3c; // 0x0a0
	13'h0a1: qq = 8'h85; // 0x0a1
	13'h0a2: qq = 8'h24; // 0x0a2
	13'h0a3: qq = 8'hbd; // 0x0a3
	13'h0a4: qq = 8'h72; // 0x0a4
	13'h0a5: qq = 8'h3c; // 0x0a5
	13'h0a6: qq = 8'h85; // 0x0a6
	13'h0a7: qq = 8'h25; // 0x0a7
	13'h0a8: qq = 8'ha0; // 0x0a8
	13'h0a9: qq = 8'h00; // 0x0a9
	13'h0aa: qq = 8'hb1; // 0x0aa
	13'h0ab: qq = 8'h22; // 0x0ab
	13'h0ac: qq = 8'hf0; // 0x0ac
	13'h0ad: qq = 8'h08; // 0x0ad
	13'h0ae: qq = 8'h05; // 0x0ae
	13'h0af: qq = 8'h28; // 0x0af
	13'h0b0: qq = 8'h91; // 0x0b0
	13'h0b1: qq = 8'h24; // 0x0b1
	13'h0b2: qq = 8'hc8; // 0x0b2
	13'h0b3: qq = 8'h4c; // 0x0b3
	13'h0b4: qq = 8'haa; // 0x0b4
	13'h0b5: qq = 8'h38; // 0x0b5
	13'h0b6: qq = 8'h60; // 0x0b6
	13'h0b7: qq = 8'hbd; // 0x0b7
	13'h0b8: qq = 8'h71; // 0x0b8
	13'h0b9: qq = 8'h3c; // 0x0b9
	13'h0ba: qq = 8'h85; // 0x0ba
	13'h0bb: qq = 8'h22; // 0x0bb
	13'h0bc: qq = 8'hbd; // 0x0bc
	13'h0bd: qq = 8'h72; // 0x0bd
	13'h0be: qq = 8'h3c; // 0x0be
	13'h0bf: qq = 8'h85; // 0x0bf
	13'h0c0: qq = 8'h23; // 0x0c0
	13'h0c1: qq = 8'ha9; // 0x0c1
	13'h0c2: qq = 8'h20; // 0x0c2
	13'h0c3: qq = 8'ha0; // 0x0c3
	13'h0c4: qq = 8'h00; // 0x0c4
	13'h0c5: qq = 8'h91; // 0x0c5
	13'h0c6: qq = 8'h22; // 0x0c6
	13'h0c7: qq = 8'hc8; // 0x0c7
	13'h0c8: qq = 8'hc0; // 0x0c8
	13'h0c9: qq = 8'h20; // 0x0c9
	13'h0ca: qq = 8'hd0; // 0x0ca
	13'h0cb: qq = 8'hf9; // 0x0cb
	13'h0cc: qq = 8'h60; // 0x0cc
	13'h0cd: qq = 8'h8d; // 0x0cd
	13'h0ce: qq = 8'h80; // 0x0ce
	13'h0cf: qq = 8'h0c; // 0x0cf
	13'h0d0: qq = 8'ha5; // 0x0d0
	13'h0d1: qq = 8'h38; // 0x0d1
	13'h0d2: qq = 8'hd0; // 0x0d2
	13'h0d3: qq = 8'h29; // 0x0d3
	13'h0d4: qq = 8'ha5; // 0x0d4
	13'h0d5: qq = 8'h35; // 0x0d5
	13'h0d6: qq = 8'hd0; // 0x0d6
	13'h0d7: qq = 8'h0d; // 0x0d7
	13'h0d8: qq = 8'ha2; // 0x0d8
	13'h0d9: qq = 8'h22; // 0x0d9
	13'h0da: qq = 8'h20; // 0x0da
	13'h0db: qq = 8'hb7; // 0x0db
	13'h0dc: qq = 8'h38; // 0x0dc
	13'h0dd: qq = 8'he8; // 0x0dd
	13'h0de: qq = 8'he8; // 0x0de
	13'h0df: qq = 8'he0; // 0x0df
	13'h0e0: qq = 8'h30; // 0x0e0
	13'h0e1: qq = 8'hd0; // 0x0e1
	13'h0e2: qq = 8'hf7; // 0x0e2
	13'h0e3: qq = 8'ha5; // 0x0e3
	13'h0e4: qq = 8'h35; // 0x0e4
	13'h0e5: qq = 8'h0a; // 0x0e5
	13'h0e6: qq = 8'haa; // 0x0e6
	13'h0e7: qq = 8'hbd; // 0x0e7
	13'h0e8: qq = 8'h37; // 0x0e8
	13'h0e9: qq = 8'h3c; // 0x0e9
	13'h0ea: qq = 8'h85; // 0x0ea
	13'h0eb: qq = 8'h24; // 0x0eb
	13'h0ec: qq = 8'hbd; // 0x0ec
	13'h0ed: qq = 8'h38; // 0x0ed
	13'h0ee: qq = 8'h3c; // 0x0ee
	13'h0ef: qq = 8'h85; // 0x0ef
	13'h0f0: qq = 8'h25; // 0x0f0
	13'h0f1: qq = 8'ha0; // 0x0f1
	13'h0f2: qq = 8'h00; // 0x0f2
	13'h0f3: qq = 8'hb1; // 0x0f3
	13'h0f4: qq = 8'h24; // 0x0f4
	13'h0f5: qq = 8'h99; // 0x0f5
	13'h0f6: qq = 8'h48; // 0x0f6
	13'h0f7: qq = 8'h00; // 0x0f7
	13'h0f8: qq = 8'hc8; // 0x0f8
	13'h0f9: qq = 8'hc0; // 0x0f9
	13'h0fa: qq = 8'h06; // 0x0fa
	13'h0fb: qq = 8'hd0; // 0x0fb
	13'h0fc: qq = 8'hf6; // 0x0fc
	13'h0fd: qq = 8'h18; // 0x0fd
	13'h0fe: qq = 8'ha5; // 0x0fe
	13'h0ff: qq = 8'h48; // 0x0ff
	13'h100: qq = 8'h69; // 0x100
	13'h101: qq = 8'h18; // 0x101
	13'h102: qq = 8'h85; // 0x102
	13'h103: qq = 8'h4e; // 0x103
	13'h104: qq = 8'ha9; // 0x104
	13'h105: qq = 8'h00; // 0x105
	13'h106: qq = 8'h65; // 0x106
	13'h107: qq = 8'h49; // 0x107
	13'h108: qq = 8'h85; // 0x108
	13'h109: qq = 8'h4f; // 0x109
	13'h10a: qq = 8'ha9; // 0x10a
	13'h10b: qq = 8'h01; // 0x10b
	13'h10c: qq = 8'h85; // 0x10c
	13'h10d: qq = 8'h38; // 0x10d
	13'h10e: qq = 8'h20; // 0x10e
	13'h10f: qq = 8'hff; // 0x10f
	13'h110: qq = 8'h37; // 0x110
	13'h111: qq = 8'ha0; // 0x111
	13'h112: qq = 8'h00; // 0x112
	13'h113: qq = 8'hb1; // 0x113
	13'h114: qq = 8'h48; // 0x114
	13'h115: qq = 8'h29; // 0x115
	13'h116: qq = 8'hf0; // 0x116
	13'h117: qq = 8'h4a; // 0x117
	13'h118: qq = 8'h4a; // 0x118
	13'h119: qq = 8'h4a; // 0x119
	13'h11a: qq = 8'h4a; // 0x11a
	13'h11b: qq = 8'h09; // 0x11b
	13'h11c: qq = 8'ha0; // 0x11c
	13'h11d: qq = 8'h91; // 0x11d
	13'h11e: qq = 8'h4c; // 0x11e
	13'h11f: qq = 8'ha5; // 0x11f
	13'h120: qq = 8'h4c; // 0x120
	13'h121: qq = 8'h18; // 0x121
	13'h122: qq = 8'h69; // 0x122
	13'h123: qq = 8'h01; // 0x123
	13'h124: qq = 8'h85; // 0x124
	13'h125: qq = 8'h4c; // 0x125
	13'h126: qq = 8'ha9; // 0x126
	13'h127: qq = 8'h00; // 0x127
	13'h128: qq = 8'h65; // 0x128
	13'h129: qq = 8'h4d; // 0x129
	13'h12a: qq = 8'h85; // 0x12a
	13'h12b: qq = 8'h4d; // 0x12b
	13'h12c: qq = 8'hb1; // 0x12c
	13'h12d: qq = 8'h48; // 0x12d
	13'h12e: qq = 8'h29; // 0x12e
	13'h12f: qq = 8'h0f; // 0x12f
	13'h130: qq = 8'h09; // 0x130
	13'h131: qq = 8'ha0; // 0x131
	13'h132: qq = 8'h91; // 0x132
	13'h133: qq = 8'h4c; // 0x133
	13'h134: qq = 8'ha5; // 0x134
	13'h135: qq = 8'h48; // 0x135
	13'h136: qq = 8'h18; // 0x136
	13'h137: qq = 8'h69; // 0x137
	13'h138: qq = 8'h01; // 0x138
	13'h139: qq = 8'h85; // 0x139
	13'h13a: qq = 8'h48; // 0x13a
	13'h13b: qq = 8'ha9; // 0x13b
	13'h13c: qq = 8'h00; // 0x13c
	13'h13d: qq = 8'h65; // 0x13d
	13'h13e: qq = 8'h49; // 0x13e
	13'h13f: qq = 8'h85; // 0x13f
	13'h140: qq = 8'h49; // 0x140
	13'h141: qq = 8'ha5; // 0x141
	13'h142: qq = 8'h4c; // 0x142
	13'h143: qq = 8'h18; // 0x143
	13'h144: qq = 8'h69; // 0x144
	13'h145: qq = 8'h01; // 0x145
	13'h146: qq = 8'h85; // 0x146
	13'h147: qq = 8'h4c; // 0x147
	13'h148: qq = 8'ha9; // 0x148
	13'h149: qq = 8'h00; // 0x149
	13'h14a: qq = 8'h65; // 0x14a
	13'h14b: qq = 8'h4d; // 0x14b
	13'h14c: qq = 8'h85; // 0x14c
	13'h14d: qq = 8'h4d; // 0x14d
	13'h14e: qq = 8'ha5; // 0x14e
	13'h14f: qq = 8'h49; // 0x14f
	13'h150: qq = 8'hc5; // 0x150
	13'h151: qq = 8'h4b; // 0x151
	13'h152: qq = 8'hf0; // 0x152
	13'h153: qq = 8'h0c; // 0x153
	13'h154: qq = 8'ha5; // 0x154
	13'h155: qq = 8'h35; // 0x155
	13'h156: qq = 8'hf0; // 0x156
	13'h157: qq = 8'hbb; // 0x157
	13'h158: qq = 8'ha5; // 0x158
	13'h159: qq = 8'h49; // 0x159
	13'h15a: qq = 8'hc5; // 0x15a
	13'h15b: qq = 8'h4f; // 0x15b
	13'h15c: qq = 8'hf0; // 0x15c
	13'h15d: qq = 8'h0e; // 0x15d
	13'h15e: qq = 8'hd0; // 0x15e
	13'h15f: qq = 8'hb3; // 0x15f
	13'h160: qq = 8'ha5; // 0x160
	13'h161: qq = 8'h48; // 0x161
	13'h162: qq = 8'hc5; // 0x162
	13'h163: qq = 8'h4a; // 0x163
	13'h164: qq = 8'hd0; // 0x164
	13'h165: qq = 8'hee; // 0x165
	13'h166: qq = 8'ha9; // 0x166
	13'h167: qq = 8'h00; // 0x167
	13'h168: qq = 8'h85; // 0x168
	13'h169: qq = 8'h38; // 0x169
	13'h16a: qq = 8'hf0; // 0x16a
	13'h16b: qq = 8'h06; // 0x16b
	13'h16c: qq = 8'ha5; // 0x16c
	13'h16d: qq = 8'h48; // 0x16d
	13'h16e: qq = 8'hc5; // 0x16e
	13'h16f: qq = 8'h4e; // 0x16f
	13'h170: qq = 8'hd0; // 0x170
	13'h171: qq = 8'ha1; // 0x171
	13'h172: qq = 8'h20; // 0x172
	13'h173: qq = 8'hff; // 0x173
	13'h174: qq = 8'h37; // 0x174
	13'h175: qq = 8'h2c; // 0x175
	13'h176: qq = 8'h30; // 0x176
	13'h177: qq = 8'h08; // 0x177
	13'h178: qq = 8'h30; // 0x178
	13'h179: qq = 8'h3c; // 0x179
	13'h17a: qq = 8'ha5; // 0x17a
	13'h17b: qq = 8'h35; // 0x17b
	13'h17c: qq = 8'h0a; // 0x17c
	13'h17d: qq = 8'h0a; // 0x17d
	13'h17e: qq = 8'ha8; // 0x17e
	13'h17f: qq = 8'ha2; // 0x17f
	13'h180: qq = 8'h00; // 0x180
	13'h181: qq = 8'hb9; // 0x181
	13'h182: qq = 8'hd6; // 0x182
	13'h183: qq = 8'h2e; // 0x183
	13'h184: qq = 8'h95; // 0x184
	13'h185: qq = 8'h22; // 0x185
	13'h186: qq = 8'hc8; // 0x186
	13'h187: qq = 8'he8; // 0x187
	13'h188: qq = 8'he0; // 0x188
	13'h189: qq = 8'h04; // 0x189
	13'h18a: qq = 8'hd0; // 0x18a
	13'h18b: qq = 8'hf5; // 0x18b
	13'h18c: qq = 8'ha2; // 0x18c
	13'h18d: qq = 8'h00; // 0x18d
	13'h18e: qq = 8'ha0; // 0x18e
	13'h18f: qq = 8'h00; // 0x18f
	13'h190: qq = 8'ha9; // 0x190
	13'h191: qq = 8'h3c; // 0x191
	13'h192: qq = 8'h91; // 0x192
	13'h193: qq = 8'h22; // 0x193
	13'h194: qq = 8'ha0; // 0x194
	13'h195: qq = 8'h01; // 0x195
	13'h196: qq = 8'ha9; // 0x196
	13'h197: qq = 8'h3d; // 0x197
	13'h198: qq = 8'h91; // 0x198
	13'h199: qq = 8'h22; // 0x199
	13'h19a: qq = 8'ha0; // 0x19a
	13'h19b: qq = 8'h20; // 0x19b
	13'h19c: qq = 8'ha9; // 0x19c
	13'h19d: qq = 8'h3e; // 0x19d
	13'h19e: qq = 8'h91; // 0x19e
	13'h19f: qq = 8'h22; // 0x19f
	13'h1a0: qq = 8'ha0; // 0x1a0
	13'h1a1: qq = 8'h21; // 0x1a1
	13'h1a2: qq = 8'ha9; // 0x1a2
	13'h1a3: qq = 8'h3f; // 0x1a3
	13'h1a4: qq = 8'h91; // 0x1a4
	13'h1a5: qq = 8'h22; // 0x1a5
	13'h1a6: qq = 8'he8; // 0x1a6
	13'h1a7: qq = 8'he0; // 0x1a7
	13'h1a8: qq = 8'h01; // 0x1a8
	13'h1a9: qq = 8'hd0; // 0x1a9
	13'h1aa: qq = 8'h0b; // 0x1aa
	13'h1ab: qq = 8'ha5; // 0x1ab
	13'h1ac: qq = 8'h24; // 0x1ac
	13'h1ad: qq = 8'h85; // 0x1ad
	13'h1ae: qq = 8'h22; // 0x1ae
	13'h1af: qq = 8'ha5; // 0x1af
	13'h1b0: qq = 8'h25; // 0x1b0
	13'h1b1: qq = 8'h85; // 0x1b1
	13'h1b2: qq = 8'h23; // 0x1b2
	13'h1b3: qq = 8'h4c; // 0x1b3
	13'h1b4: qq = 8'h8e; // 0x1b4
	13'h1b5: qq = 8'h39; // 0x1b5
	13'h1b6: qq = 8'h8d; // 0x1b6
	13'h1b7: qq = 8'h80; // 0x1b7
	13'h1b8: qq = 8'h0c; // 0x1b8
	13'h1b9: qq = 8'h60; // 0x1b9
	13'h1ba: qq = 8'had; // 0x1ba
	13'h1bb: qq = 8'h6b; // 0x1bb
	13'h1bc: qq = 8'h04; // 0x1bc
	13'h1bd: qq = 8'hc9; // 0x1bd
	13'h1be: qq = 8'hcb; // 0x1be
	13'h1bf: qq = 8'hd0; // 0x1bf
	13'h1c0: qq = 8'h26; // 0x1c0
	13'h1c1: qq = 8'had; // 0x1c1
	13'h1c2: qq = 8'h04; // 0x1c2
	13'h1c3: qq = 8'h3e; // 0x1c3
	13'h1c4: qq = 8'hc9; // 0x1c4
	13'h1c5: qq = 8'h4b; // 0x1c5
	13'h1c6: qq = 8'hd0; // 0x1c6
	13'h1c7: qq = 8'h1f; // 0x1c7
	13'h1c8: qq = 8'h2c; // 0x1c8
	13'h1c9: qq = 8'h2f; // 0x1c9
	13'h1ca: qq = 8'h08; // 0x1ca
	13'h1cb: qq = 8'h30; // 0x1cb
	13'h1cc: qq = 8'h01; // 0x1cc
	13'h1cd: qq = 8'h60; // 0x1cd
	13'h1ce: qq = 8'h2c; // 0x1ce
	13'h1cf: qq = 8'h00; // 0x1cf
	13'h1d0: qq = 8'h0c; // 0x1d0
	13'h1d1: qq = 8'h10; // 0x1d1
	13'h1d2: qq = 8'hfb; // 0x1d2
	13'h1d3: qq = 8'h2c; // 0x1d3
	13'h1d4: qq = 8'h00; // 0x1d4
	13'h1d5: qq = 8'h0c; // 0x1d5
	13'h1d6: qq = 8'h30; // 0x1d6
	13'h1d7: qq = 8'hfb; // 0x1d7
	13'h1d8: qq = 8'ha9; // 0x1d8
	13'h1d9: qq = 8'h0a; // 0x1d9
	13'h1da: qq = 8'ha0; // 0x1da
	13'h1db: qq = 8'h00; // 0x1db
	13'h1dc: qq = 8'hc8; // 0x1dc
	13'h1dd: qq = 8'hd0; // 0x1dd
	13'h1de: qq = 8'hfd; // 0x1de
	13'h1df: qq = 8'h38; // 0x1df
	13'h1e0: qq = 8'he9; // 0x1e0
	13'h1e1: qq = 8'h01; // 0x1e1
	13'h1e2: qq = 8'hd0; // 0x1e2
	13'h1e3: qq = 8'hf6; // 0x1e3
	13'h1e4: qq = 8'h30; // 0x1e4
	13'h1e5: qq = 8'h01; // 0x1e5
	13'h1e6: qq = 8'h60; // 0x1e6
	13'h1e7: qq = 8'ha9; // 0x1e7
	13'h1e8: qq = 8'h00; // 0x1e8
	13'h1e9: qq = 8'h85; // 0x1e9
	13'h1ea: qq = 8'h20; // 0x1ea
	13'h1eb: qq = 8'h85; // 0x1eb
	13'h1ec: qq = 8'h36; // 0x1ec
	13'h1ed: qq = 8'h60; // 0x1ed
	13'h1ee: qq = 8'ha9; // 0x1ee
	13'h1ef: qq = 8'h00; // 0x1ef
	13'h1f0: qq = 8'ha2; // 0x1f0
	13'h1f1: qq = 8'h20; // 0x1f1
	13'h1f2: qq = 8'h20; // 0x1f2
	13'h1f3: qq = 8'h8a; // 0x1f3
	13'h1f4: qq = 8'h38; // 0x1f4
	13'h1f5: qq = 8'had; // 0x1f5
	13'h1f6: qq = 8'h28; // 0x1f6
	13'h1f7: qq = 8'h04; // 0x1f7
	13'h1f8: qq = 8'h29; // 0x1f8
	13'h1f9: qq = 8'h3f; // 0x1f9
	13'h1fa: qq = 8'hc5; // 0x1fa
	13'h1fb: qq = 8'h59; // 0x1fb
	13'h1fc: qq = 8'h30; // 0x1fc
	13'h1fd: qq = 8'h2f; // 0x1fd
	13'h1fe: qq = 8'hf0; // 0x1fe
	13'h1ff: qq = 8'h02; // 0x1ff
	13'h200: qq = 8'h10; // 0x200
	13'h201: qq = 8'h16; // 0x201
	13'h202: qq = 8'had; // 0x202
	13'h203: qq = 8'h29; // 0x203
	13'h204: qq = 8'h04; // 0x204
	13'h205: qq = 8'h29; // 0x205
	13'h206: qq = 8'h3f; // 0x206
	13'h207: qq = 8'hc5; // 0x207
	13'h208: qq = 8'h58; // 0x208
	13'h209: qq = 8'h30; // 0x209
	13'h20a: qq = 8'h22; // 0x20a
	13'h20b: qq = 8'hf0; // 0x20b
	13'h20c: qq = 8'h02; // 0x20c
	13'h20d: qq = 8'h10; // 0x20d
	13'h20e: qq = 8'h09; // 0x20e
	13'h20f: qq = 8'had; // 0x20f
	13'h210: qq = 8'h2a; // 0x210
	13'h211: qq = 8'h04; // 0x211
	13'h212: qq = 8'h29; // 0x212
	13'h213: qq = 8'h3f; // 0x213
	13'h214: qq = 8'hc5; // 0x214
	13'h215: qq = 8'h57; // 0x215
	13'h216: qq = 8'h30; // 0x216
	13'h217: qq = 8'h15; // 0x217
	13'h218: qq = 8'had; // 0x218
	13'h219: qq = 8'h28; // 0x219
	13'h21a: qq = 8'h04; // 0x21a
	13'h21b: qq = 8'h29; // 0x21b
	13'h21c: qq = 8'h3f; // 0x21c
	13'h21d: qq = 8'h85; // 0x21d
	13'h21e: qq = 8'h59; // 0x21e
	13'h21f: qq = 8'had; // 0x21f
	13'h220: qq = 8'h29; // 0x220
	13'h221: qq = 8'h04; // 0x221
	13'h222: qq = 8'h29; // 0x222
	13'h223: qq = 8'h3f; // 0x223
	13'h224: qq = 8'h85; // 0x224
	13'h225: qq = 8'h58; // 0x225
	13'h226: qq = 8'had; // 0x226
	13'h227: qq = 8'h2a; // 0x227
	13'h228: qq = 8'h04; // 0x228
	13'h229: qq = 8'h29; // 0x229
	13'h22a: qq = 8'h3f; // 0x22a
	13'h22b: qq = 8'h85; // 0x22b
	13'h22c: qq = 8'h57; // 0x22c
	13'h22d: qq = 8'ha5; // 0x22d
	13'h22e: qq = 8'h57; // 0x22e
	13'h22f: qq = 8'h8d; // 0x22f
	13'h230: qq = 8'h3b; // 0x230
	13'h231: qq = 8'h04; // 0x231
	13'h232: qq = 8'ha5; // 0x232
	13'h233: qq = 8'h58; // 0x233
	13'h234: qq = 8'h8d; // 0x234
	13'h235: qq = 8'h3a; // 0x235
	13'h236: qq = 8'h04; // 0x236
	13'h237: qq = 8'ha5; // 0x237
	13'h238: qq = 8'h59; // 0x238
	13'h239: qq = 8'h8d; // 0x239
	13'h23a: qq = 8'h39; // 0x23a
	13'h23b: qq = 8'h04; // 0x23b
	13'h23c: qq = 8'h60; // 0x23c
	13'h23d: qq = 8'ha2; // 0x23d
	13'h23e: qq = 8'h00; // 0x23e
	13'h23f: qq = 8'ha0; // 0x23f
	13'h240: qq = 8'h00; // 0x240
	13'h241: qq = 8'hb5; // 0x241
	13'h242: qq = 8'h40; // 0x242
	13'h243: qq = 8'h95; // 0x243
	13'h244: qq = 8'h10; // 0x244
	13'h245: qq = 8'hb5; // 0x245
	13'h246: qq = 8'h44; // 0x246
	13'h247: qq = 8'h99; // 0x247
	13'h248: qq = 8'h18; // 0x248
	13'h249: qq = 8'h00; // 0x249
	13'h24a: qq = 8'he8; // 0x24a
	13'h24b: qq = 8'hc8; // 0x24b
	13'h24c: qq = 8'hc8; // 0x24c
	13'h24d: qq = 8'he0; // 0x24d
	13'h24e: qq = 8'h04; // 0x24e
	13'h24f: qq = 8'hd0; // 0x24f
	13'h250: qq = 8'hf0; // 0x250
	13'h251: qq = 8'h60; // 0x251
	13'h252: qq = 8'ha2; // 0x252
	13'h253: qq = 8'h00; // 0x253
	13'h254: qq = 8'ha9; // 0x254
	13'h255: qq = 8'h01; // 0x255
	13'h256: qq = 8'h9d; // 0x256
	13'h257: qq = 8'h00; // 0x257
	13'h258: qq = 8'h04; // 0x258
	13'h259: qq = 8'h8d; // 0x259
	13'h25a: qq = 8'h80; // 0x25a
	13'h25b: qq = 8'h0c; // 0x25b
	13'h25c: qq = 8'hdd; // 0x25c
	13'h25d: qq = 8'h00; // 0x25d
	13'h25e: qq = 8'h04; // 0x25e
	13'h25f: qq = 8'hd0; // 0x25f
	13'h260: qq = 8'hf5; // 0x260
	13'h261: qq = 8'h9d; // 0x261
	13'h262: qq = 8'h00; // 0x262
	13'h263: qq = 8'h05; // 0x263
	13'h264: qq = 8'h8d; // 0x264
	13'h265: qq = 8'h80; // 0x265
	13'h266: qq = 8'h0c; // 0x266
	13'h267: qq = 8'hdd; // 0x267
	13'h268: qq = 8'h00; // 0x268
	13'h269: qq = 8'h05; // 0x269
	13'h26a: qq = 8'hd0; // 0x26a
	13'h26b: qq = 8'hf5; // 0x26b
	13'h26c: qq = 8'h9d; // 0x26c
	13'h26d: qq = 8'h00; // 0x26d
	13'h26e: qq = 8'h06; // 0x26e
	13'h26f: qq = 8'h8d; // 0x26f
	13'h270: qq = 8'h80; // 0x270
	13'h271: qq = 8'h0c; // 0x271
	13'h272: qq = 8'hdd; // 0x272
	13'h273: qq = 8'h00; // 0x273
	13'h274: qq = 8'h06; // 0x274
	13'h275: qq = 8'hd0; // 0x275
	13'h276: qq = 8'hf5; // 0x276
	13'h277: qq = 8'h9d; // 0x277
	13'h278: qq = 8'h00; // 0x278
	13'h279: qq = 8'h07; // 0x279
	13'h27a: qq = 8'h8d; // 0x27a
	13'h27b: qq = 8'h80; // 0x27b
	13'h27c: qq = 8'h0c; // 0x27c
	13'h27d: qq = 8'hdd; // 0x27d
	13'h27e: qq = 8'h00; // 0x27e
	13'h27f: qq = 8'h07; // 0x27f
	13'h280: qq = 8'hd0; // 0x280
	13'h281: qq = 8'hf5; // 0x281
	13'h282: qq = 8'he8; // 0x282
	13'h283: qq = 8'hd0; // 0x283
	13'h284: qq = 8'hd1; // 0x284
	13'h285: qq = 8'h18; // 0x285
	13'h286: qq = 8'h69; // 0x286
	13'h287: qq = 8'h01; // 0x287
	13'h288: qq = 8'hc9; // 0x288
	13'h289: qq = 8'h01; // 0x289
	13'h28a: qq = 8'hd0; // 0x28a
	13'h28b: qq = 8'hca; // 0x28b
	13'h28c: qq = 8'ha9; // 0x28c
	13'h28d: qq = 8'h00; // 0x28d
	13'h28e: qq = 8'h85; // 0x28e
	13'h28f: qq = 8'h16; // 0x28f
	13'h290: qq = 8'ha2; // 0x290
	13'h291: qq = 8'h00; // 0x291
	13'h292: qq = 8'ha9; // 0x292
	13'h293: qq = 8'h10; // 0x293
	13'h294: qq = 8'h85; // 0x294
	13'h295: qq = 8'h24; // 0x295
	13'h296: qq = 8'ha9; // 0x296
	13'h297: qq = 8'h05; // 0x297
	13'h298: qq = 8'h85; // 0x298
	13'h299: qq = 8'h25; // 0x299
	13'h29a: qq = 8'ha9; // 0x29a
	13'h29b: qq = 8'h00; // 0x29b
	13'h29c: qq = 8'h85; // 0x29c
	13'h29d: qq = 8'h7e; // 0x29d
	13'h29e: qq = 8'ha9; // 0x29e
	13'h29f: qq = 8'h20; // 0x29f
	13'h2a0: qq = 8'h85; // 0x2a0
	13'h2a1: qq = 8'h7f; // 0x2a1
	13'h2a2: qq = 8'ha0; // 0x2a2
	13'h2a3: qq = 8'h00; // 0x2a3
	13'h2a4: qq = 8'ha9; // 0x2a4
	13'h2a5: qq = 8'h00; // 0x2a5
	13'h2a6: qq = 8'h85; // 0x2a6
	13'h2a7: qq = 8'h26; // 0x2a7
	13'h2a8: qq = 8'h85; // 0x2a8
	13'h2a9: qq = 8'h22; // 0x2a9
	13'h2aa: qq = 8'ha5; // 0x2aa
	13'h2ab: qq = 8'h22; // 0x2ab
	13'h2ac: qq = 8'h18; // 0x2ac
	13'h2ad: qq = 8'h71; // 0x2ad
	13'h2ae: qq = 8'h7e; // 0x2ae
	13'h2af: qq = 8'h85; // 0x2af
	13'h2b0: qq = 8'h22; // 0x2b0
	13'h2b1: qq = 8'hc8; // 0x2b1
	13'h2b2: qq = 8'hd0; // 0x2b2
	13'h2b3: qq = 8'hf6; // 0x2b3
	13'h2b4: qq = 8'h8d; // 0x2b4
	13'h2b5: qq = 8'h80; // 0x2b5
	13'h2b6: qq = 8'h0c; // 0x2b6
	13'h2b7: qq = 8'he6; // 0x2b7
	13'h2b8: qq = 8'h7f; // 0x2b8
	13'h2b9: qq = 8'he6; // 0x2b9
	13'h2ba: qq = 8'h26; // 0x2ba
	13'h2bb: qq = 8'ha5; // 0x2bb
	13'h2bc: qq = 8'h26; // 0x2bc
	13'h2bd: qq = 8'hc9; // 0x2bd
	13'h2be: qq = 8'h04; // 0x2be
	13'h2bf: qq = 8'hd0; // 0x2bf
	13'h2c0: qq = 8'he9; // 0x2c0
	13'h2c1: qq = 8'ha5; // 0x2c1
	13'h2c2: qq = 8'h22; // 0x2c2
	13'h2c3: qq = 8'hdd; // 0x2c3
	13'h2c4: qq = 8'h2e; // 0x2c4
	13'h2c5: qq = 8'h3c; // 0x2c5
	13'h2c6: qq = 8'hf0; // 0x2c6
	13'h2c7: qq = 8'h09; // 0x2c7
	13'h2c8: qq = 8'ha0; // 0x2c8
	13'h2c9: qq = 8'h00; // 0x2c9
	13'h2ca: qq = 8'h8a; // 0x2ca
	13'h2cb: qq = 8'h09; // 0x2cb
	13'h2cc: qq = 8'h30; // 0x2cc
	13'h2cd: qq = 8'h91; // 0x2cd
	13'h2ce: qq = 8'h24; // 0x2ce
	13'h2cf: qq = 8'he6; // 0x2cf
	13'h2d0: qq = 8'h24; // 0x2d0
	13'h2d1: qq = 8'he8; // 0x2d1
	13'h2d2: qq = 8'he0; // 0x2d2
	13'h2d3: qq = 8'h08; // 0x2d3
	13'h2d4: qq = 8'hd0; // 0x2d4
	13'h2d5: qq = 8'hcc; // 0x2d5
	13'h2d6: qq = 8'ha9; // 0x2d6
	13'h2d7: qq = 8'hd4; // 0x2d7
	13'h2d8: qq = 8'h8d; // 0x2d8
	13'h2d9: qq = 8'h6a; // 0x2d9
	13'h2da: qq = 8'h04; // 0x2da
	13'h2db: qq = 8'ha9; // 0x2db
	13'h2dc: qq = 8'hc9; // 0x2dc
	13'h2dd: qq = 8'h8d; // 0x2dd
	13'h2de: qq = 8'h6b; // 0x2de
	13'h2df: qq = 8'h04; // 0x2df
	13'h2e0: qq = 8'ha9; // 0x2e0
	13'h2e1: qq = 8'hcd; // 0x2e1
	13'h2e2: qq = 8'h8d; // 0x2e2
	13'h2e3: qq = 8'h6c; // 0x2e3
	13'h2e4: qq = 8'h04; // 0x2e4
	13'h2e5: qq = 8'ha9; // 0x2e5
	13'h2e6: qq = 8'hc5; // 0x2e6
	13'h2e7: qq = 8'h8d; // 0x2e7
	13'h2e8: qq = 8'h6d; // 0x2e8
	13'h2e9: qq = 8'h04; // 0x2e9
	13'h2ea: qq = 8'ha9; // 0x2ea
	13'h2eb: qq = 8'hcc; // 0x2eb
	13'h2ec: qq = 8'h8d; // 0x2ec
	13'h2ed: qq = 8'hcc; // 0x2ed
	13'h2ee: qq = 8'h04; // 0x2ee
	13'h2ef: qq = 8'ha9; // 0x2ef
	13'h2f0: qq = 8'hc1; // 0x2f0
	13'h2f1: qq = 8'h8d; // 0x2f1
	13'h2f2: qq = 8'hcd; // 0x2f2
	13'h2f3: qq = 8'h04; // 0x2f3
	13'h2f4: qq = 8'ha9; // 0x2f4
	13'h2f5: qq = 8'hd0; // 0x2f5
	13'h2f6: qq = 8'h8d; // 0x2f6
	13'h2f7: qq = 8'hce; // 0x2f7
	13'h2f8: qq = 8'h04; // 0x2f8
	13'h2f9: qq = 8'ha9; // 0x2f9
	13'h2fa: qq = 8'hd3; // 0x2fa
	13'h2fb: qq = 8'h8d; // 0x2fb
	13'h2fc: qq = 8'hcf; // 0x2fc
	13'h2fd: qq = 8'h04; // 0x2fd
	13'h2fe: qq = 8'ha9; // 0x2fe
	13'h2ff: qq = 8'hb0; // 0x2ff
	13'h300: qq = 8'h8d; // 0x300
	13'h301: qq = 8'h71; // 0x301
	13'h302: qq = 8'h04; // 0x302
	13'h303: qq = 8'ha9; // 0x303
	13'h304: qq = 8'hb1; // 0x304
	13'h305: qq = 8'h2c; // 0x305
	13'h306: qq = 8'h30; // 0x306
	13'h307: qq = 8'h08; // 0x307
	13'h308: qq = 8'h70; // 0x308
	13'h309: qq = 8'h02; // 0x309
	13'h30a: qq = 8'ha9; // 0x30a
	13'h30b: qq = 8'hb2; // 0x30b
	13'h30c: qq = 8'h8d; // 0x30c
	13'h30d: qq = 8'hca; // 0x30d
	13'h30e: qq = 8'h04; // 0x30e
	13'h30f: qq = 8'ha9; // 0x30f
	13'h310: qq = 8'h20; // 0x310
	13'h311: qq = 8'h2c; // 0x311
	13'h312: qq = 8'h33; // 0x312
	13'h313: qq = 8'h08; // 0x313
	13'h314: qq = 8'h30; // 0x314
	13'h315: qq = 8'h02; // 0x315
	13'h316: qq = 8'ha9; // 0x316
	13'h317: qq = 8'hb1; // 0x317
	13'h318: qq = 8'h8d; // 0x318
	13'h319: qq = 8'h6f; // 0x319
	13'h31a: qq = 8'h04; // 0x31a
	13'h31b: qq = 8'ha9; // 0x31b
	13'h31c: qq = 8'hb6; // 0x31c
	13'h31d: qq = 8'h2c; // 0x31d
	13'h31e: qq = 8'h33; // 0x31e
	13'h31f: qq = 8'h08; // 0x31f
	13'h320: qq = 8'h30; // 0x320
	13'h321: qq = 8'h08; // 0x321
	13'h322: qq = 8'ha9; // 0x322
	13'h323: qq = 8'hb2; // 0x323
	13'h324: qq = 8'h70; // 0x324
	13'h325: qq = 8'h02; // 0x325
	13'h326: qq = 8'ha9; // 0x326
	13'h327: qq = 8'hb5; // 0x327
	13'h328: qq = 8'h30; // 0x328
	13'h329: qq = 8'h04; // 0x329
	13'h32a: qq = 8'h70; // 0x32a
	13'h32b: qq = 8'h02; // 0x32b
	13'h32c: qq = 8'ha9; // 0x32c
	13'h32d: qq = 8'hb9; // 0x32d
	13'h32e: qq = 8'h8d; // 0x32e
	13'h32f: qq = 8'h70; // 0x32f
	13'h330: qq = 8'h04; // 0x330
	13'h331: qq = 8'ha9; // 0x331
	13'h332: qq = 8'h8a; // 0x332
	13'h333: qq = 8'h85; // 0x333
	13'h334: qq = 8'h22; // 0x334
	13'h335: qq = 8'ha9; // 0x335
	13'h336: qq = 8'h04; // 0x336
	13'h337: qq = 8'h85; // 0x337
	13'h338: qq = 8'h23; // 0x338
	13'h339: qq = 8'h2c; // 0x339
	13'h33a: qq = 8'h31; // 0x33a
	13'h33b: qq = 8'h08; // 0x33b
	13'h33c: qq = 8'h30; // 0x33c
	13'h33d: qq = 8'h18; // 0x33d
	13'h33e: qq = 8'h70; // 0x33e
	13'h33f: qq = 8'h0b; // 0x33f
	13'h340: qq = 8'ha9; // 0x340
	13'h341: qq = 8'h05; // 0x341
	13'h342: qq = 8'h85; // 0x342
	13'h343: qq = 8'h24; // 0x343
	13'h344: qq = 8'ha9; // 0x344
	13'h345: qq = 8'h3d; // 0x345
	13'h346: qq = 8'h85; // 0x346
	13'h347: qq = 8'h25; // 0x347
	13'h348: qq = 8'h4c; // 0x348
	13'h349: qq = 8'h86; // 0x349
	13'h34a: qq = 8'h3b; // 0x34a
	13'h34b: qq = 8'ha9; // 0x34b
	13'h34c: qq = 8'h3c; // 0x34c
	13'h34d: qq = 8'h85; // 0x34d
	13'h34e: qq = 8'h24; // 0x34e
	13'h34f: qq = 8'ha9; // 0x34f
	13'h350: qq = 8'h3d; // 0x350
	13'h351: qq = 8'h85; // 0x351
	13'h352: qq = 8'h25; // 0x352
	13'h353: qq = 8'h4c; // 0x353
	13'h354: qq = 8'h86; // 0x354
	13'h355: qq = 8'h3b; // 0x355
	13'h356: qq = 8'h70; // 0x356
	13'h357: qq = 8'h0b; // 0x357
	13'h358: qq = 8'ha9; // 0x358
	13'h359: qq = 8'h20; // 0x359
	13'h35a: qq = 8'h85; // 0x35a
	13'h35b: qq = 8'h24; // 0x35b
	13'h35c: qq = 8'ha9; // 0x35c
	13'h35d: qq = 8'h3d; // 0x35d
	13'h35e: qq = 8'h85; // 0x35e
	13'h35f: qq = 8'h25; // 0x35f
	13'h360: qq = 8'h4c; // 0x360
	13'h361: qq = 8'h86; // 0x361
	13'h362: qq = 8'h3b; // 0x362
	13'h363: qq = 8'ha9; // 0x363
	13'h364: qq = 8'hc4; // 0x364
	13'h365: qq = 8'h8d; // 0x365
	13'h366: qq = 8'h8a; // 0x366
	13'h367: qq = 8'h04; // 0x367
	13'h368: qq = 8'ha9; // 0x368
	13'h369: qq = 8'hc5; // 0x369
	13'h36a: qq = 8'h8d; // 0x36a
	13'h36b: qq = 8'h8b; // 0x36b
	13'h36c: qq = 8'h04; // 0x36c
	13'h36d: qq = 8'ha9; // 0x36d
	13'h36e: qq = 8'hcd; // 0x36e
	13'h36f: qq = 8'h8d; // 0x36f
	13'h370: qq = 8'h8c; // 0x370
	13'h371: qq = 8'h04; // 0x371
	13'h372: qq = 8'ha9; // 0x372
	13'h373: qq = 8'hcf; // 0x373
	13'h374: qq = 8'h8d; // 0x374
	13'h375: qq = 8'h8d; // 0x375
	13'h376: qq = 8'h04; // 0x376
	13'h377: qq = 8'ha2; // 0x377
	13'h378: qq = 8'h00; // 0x378
	13'h379: qq = 8'ha9; // 0x379
	13'h37a: qq = 8'h20; // 0x37a
	13'h37b: qq = 8'h9d; // 0x37b
	13'h37c: qq = 8'h8e; // 0x37c
	13'h37d: qq = 8'h04; // 0x37d
	13'h37e: qq = 8'he8; // 0x37e
	13'h37f: qq = 8'he0; // 0x37f
	13'h380: qq = 8'h0c; // 0x380
	13'h381: qq = 8'hd0; // 0x381
	13'h382: qq = 8'hf8; // 0x382
	13'h383: qq = 8'h4c; // 0x383
	13'h384: qq = 8'h93; // 0x384
	13'h385: qq = 8'h3b; // 0x385
	13'h386: qq = 8'ha0; // 0x386
	13'h387: qq = 8'h00; // 0x387
	13'h388: qq = 8'hb1; // 0x388
	13'h389: qq = 8'h24; // 0x389
	13'h38a: qq = 8'h09; // 0x38a
	13'h38b: qq = 8'h80; // 0x38b
	13'h38c: qq = 8'h91; // 0x38c
	13'h38d: qq = 8'h22; // 0x38d
	13'h38e: qq = 8'hc8; // 0x38e
	13'h38f: qq = 8'hc0; // 0x38f
	13'h390: qq = 8'h10; // 0x390
	13'h391: qq = 8'hd0; // 0x391
	13'h392: qq = 8'hf5; // 0x392
	13'h393: qq = 8'h2c; // 0x393
	13'h394: qq = 8'h32; // 0x394
	13'h395: qq = 8'h08; // 0x395
	13'h396: qq = 8'h10; // 0x396
	13'h397: qq = 8'h0f; // 0x397
	13'h398: qq = 8'ha2; // 0x398
	13'h399: qq = 8'h00; // 0x399
	13'h39a: qq = 8'ha9; // 0x39a
	13'h39b: qq = 8'h20; // 0x39b
	13'h39c: qq = 8'h9d; // 0x39c
	13'h39d: qq = 8'haa; // 0x39d
	13'h39e: qq = 8'h04; // 0x39e
	13'h39f: qq = 8'he8; // 0x39f
	13'h3a0: qq = 8'he0; // 0x3a0
	13'h3a1: qq = 8'h0d; // 0x3a1
	13'h3a2: qq = 8'hd0; // 0x3a2
	13'h3a3: qq = 8'hf8; // 0x3a3
	13'h3a4: qq = 8'h4c; // 0x3a4
	13'h3a5: qq = 8'hc4; // 0x3a5
	13'h3a6: qq = 8'h3b; // 0x3a6
	13'h3a7: qq = 8'ha9; // 0x3a7
	13'h3a8: qq = 8'haa; // 0x3a8
	13'h3a9: qq = 8'h85; // 0x3a9
	13'h3aa: qq = 8'h22; // 0x3aa
	13'h3ab: qq = 8'ha9; // 0x3ab
	13'h3ac: qq = 8'h04; // 0x3ac
	13'h3ad: qq = 8'h85; // 0x3ad
	13'h3ae: qq = 8'h23; // 0x3ae
	13'h3af: qq = 8'ha9; // 0x3af
	13'h3b0: qq = 8'hd5; // 0x3b0
	13'h3b1: qq = 8'h85; // 0x3b1
	13'h3b2: qq = 8'h24; // 0x3b2
	13'h3b3: qq = 8'ha9; // 0x3b3
	13'h3b4: qq = 8'h3c; // 0x3b4
	13'h3b5: qq = 8'h85; // 0x3b5
	13'h3b6: qq = 8'h25; // 0x3b6
	13'h3b7: qq = 8'ha0; // 0x3b7
	13'h3b8: qq = 8'h00; // 0x3b8
	13'h3b9: qq = 8'hb1; // 0x3b9
	13'h3ba: qq = 8'h24; // 0x3ba
	13'h3bb: qq = 8'h09; // 0x3bb
	13'h3bc: qq = 8'h80; // 0x3bc
	13'h3bd: qq = 8'h91; // 0x3bd
	13'h3be: qq = 8'h22; // 0x3be
	13'h3bf: qq = 8'hc8; // 0x3bf
	13'h3c0: qq = 8'hc0; // 0x3c0
	13'h3c1: qq = 8'h0d; // 0x3c1
	13'h3c2: qq = 8'hd0; // 0x3c2
	13'h3c3: qq = 8'hf5; // 0x3c3
	13'h3c4: qq = 8'ha9; // 0x3c4
	13'h3c5: qq = 8'h20; // 0x3c5
	13'h3c6: qq = 8'h2c; // 0x3c6
	13'h3c7: qq = 8'h30; // 0x3c7
	13'h3c8: qq = 8'h08; // 0x3c8
	13'h3c9: qq = 8'h30; // 0x3c9
	13'h3ca: qq = 8'h02; // 0x3ca
	13'h3cb: qq = 8'ha9; // 0x3cb
	13'h3cc: qq = 8'h3c; // 0x3cc
	13'h3cd: qq = 8'h8d; // 0x3cd
	13'h3ce: qq = 8'hea; // 0x3ce
	13'h3cf: qq = 8'h04; // 0x3cf
	13'h3d0: qq = 8'h2c; // 0x3d0
	13'h3d1: qq = 8'h30; // 0x3d1
	13'h3d2: qq = 8'h08; // 0x3d2
	13'h3d3: qq = 8'h30; // 0x3d3
	13'h3d4: qq = 8'h02; // 0x3d4
	13'h3d5: qq = 8'ha9; // 0x3d5
	13'h3d6: qq = 8'h3d; // 0x3d6
	13'h3d7: qq = 8'h8d; // 0x3d7
	13'h3d8: qq = 8'heb; // 0x3d8
	13'h3d9: qq = 8'h04; // 0x3d9
	13'h3da: qq = 8'h2c; // 0x3da
	13'h3db: qq = 8'h30; // 0x3db
	13'h3dc: qq = 8'h08; // 0x3dc
	13'h3dd: qq = 8'h30; // 0x3dd
	13'h3de: qq = 8'h02; // 0x3de
	13'h3df: qq = 8'ha9; // 0x3df
	13'h3e0: qq = 8'h3e; // 0x3e0
	13'h3e1: qq = 8'h8d; // 0x3e1
	13'h3e2: qq = 8'h0a; // 0x3e2
	13'h3e3: qq = 8'h05; // 0x3e3
	13'h3e4: qq = 8'h2c; // 0x3e4
	13'h3e5: qq = 8'h30; // 0x3e5
	13'h3e6: qq = 8'h08; // 0x3e6
	13'h3e7: qq = 8'h30; // 0x3e7
	13'h3e8: qq = 8'h02; // 0x3e8
	13'h3e9: qq = 8'ha9; // 0x3e9
	13'h3ea: qq = 8'h3f; // 0x3ea
	13'h3eb: qq = 8'h8d; // 0x3eb
	13'h3ec: qq = 8'h0b; // 0x3ec
	13'h3ed: qq = 8'h05; // 0x3ed
	13'h3ee: qq = 8'h2c; // 0x3ee
	13'h3ef: qq = 8'h2c; // 0x3ef
	13'h3f0: qq = 8'h08; // 0x3f0
	13'h3f1: qq = 8'h10; // 0x3f1
	13'h3f2: qq = 8'h03; // 0x3f2
	13'h3f3: qq = 8'h4c; // 0x3f3
	13'h3f4: qq = 8'h3c; // 0x3f4
	13'h3f5: qq = 8'h30; // 0x3f5
	13'h3f6: qq = 8'h8d; // 0x3f6
	13'h3f7: qq = 8'h30; // 0x3f7
	13'h3f8: qq = 8'h0c; // 0x3f8
	13'h3f9: qq = 8'h8d; // 0x3f9
	13'h3fa: qq = 8'h10; // 0x3fa
	13'h3fb: qq = 8'h0c; // 0x3fb
	13'h3fc: qq = 8'ha2; // 0x3fc
	13'h3fd: qq = 8'h00; // 0x3fd
	13'h3fe: qq = 8'hbd; // 0x3fe
	13'h3ff: qq = 8'h28; // 0x3ff
	13'h400: qq = 8'h08; // 0x400
	13'h401: qq = 8'h8d; // 0x401
	13'h402: qq = 8'h80; // 0x402
	13'h403: qq = 8'h0c; // 0x403
	13'h404: qq = 8'h30; // 0x404
	13'h405: qq = 8'h03; // 0x405
	13'h406: qq = 8'h8d; // 0x406
	13'h407: qq = 8'h11; // 0x407
	13'h408: qq = 8'h0c; // 0x408
	13'h409: qq = 8'he8; // 0x409
	13'h40a: qq = 8'he0; // 0x40a
	13'h40b: qq = 8'h03; // 0x40b
	13'h40c: qq = 8'hd0; // 0x40c
	13'h40d: qq = 8'hf0; // 0x40d
	13'h40e: qq = 8'had; // 0x40e
	13'h40f: qq = 8'h2b; // 0x40f
	13'h410: qq = 8'h08; // 0x410
	13'h411: qq = 8'h30; // 0x411
	13'h412: qq = 8'h03; // 0x412
	13'h413: qq = 8'h8d; // 0x413
	13'h414: qq = 8'h11; // 0x414
	13'h415: qq = 8'h0c; // 0x415
	13'h416: qq = 8'h2c; // 0x416
	13'h417: qq = 8'h40; // 0x417
	13'h418: qq = 8'h08; // 0x418
	13'h419: qq = 8'h30; // 0x419
	13'h41a: qq = 8'h03; // 0x41a
	13'h41b: qq = 8'h8d; // 0x41b
	13'h41c: qq = 8'h11; // 0x41c
	13'h41d: qq = 8'h0c; // 0x41d
	13'h41e: qq = 8'h70; // 0x41e
	13'h41f: qq = 8'h03; // 0x41f
	13'h420: qq = 8'h8d; // 0x420
	13'h421: qq = 8'h11; // 0x421
	13'h422: qq = 8'h0c; // 0x422
	13'h423: qq = 8'h2c; // 0x423
	13'h424: qq = 8'h2d; // 0x424
	13'h425: qq = 8'h08; // 0x425
	13'h426: qq = 8'h30; // 0x426
	13'h427: qq = 8'h03; // 0x427
	13'h428: qq = 8'h8d; // 0x428
	13'h429: qq = 8'h11; // 0x429
	13'h42a: qq = 8'h0c; // 0x42a
	13'h42b: qq = 8'h4c; // 0x42b
	13'h42c: qq = 8'h03; // 0x42c
	13'h42d: qq = 8'h3b; // 0x42d
	13'h42e: qq = 8'hcc; // 0x42e
	13'h42f: qq = 8'h51; // 0x42f
	13'h430: qq = 8'h09; // 0x430
	13'h431: qq = 8'h91; // 0x431
	13'h432: qq = 8'h38; // 0x432
	13'h433: qq = 8'h2f; // 0x433
	13'h434: qq = 8'hac; // 0x434
	13'h435: qq = 8'h46; // 0x435
	13'h436: qq = 8'h30; // 0x436
	13'h437: qq = 8'h00; // 0x437
	13'h438: qq = 8'h20; // 0x438
	13'h439: qq = 8'h26; // 0x439
	13'h43a: qq = 8'h21; // 0x43a
	13'h43b: qq = 8'h4c; // 0x43b
	13'h43c: qq = 8'h22; // 0x43c
	13'h43d: qq = 8'h72; // 0x43d
	13'h43e: qq = 8'h23; // 0x43e
	13'h43f: qq = 8'h98; // 0x43f
	13'h440: qq = 8'h24; // 0x440
	13'h441: qq = 8'hbe; // 0x441
	13'h442: qq = 8'h25; // 0x442
	13'h443: qq = 8'he4; // 0x443
	13'h444: qq = 8'h26; // 0x444
	13'h445: qq = 8'h0a; // 0x445
	13'h446: qq = 8'h28; // 0x446
	13'h447: qq = 8'h30; // 0x447
	13'h448: qq = 8'h29; // 0x448
	13'h449: qq = 8'h56; // 0x449
	13'h44a: qq = 8'h2a; // 0x44a
	13'h44b: qq = 8'h7c; // 0x44b
	13'h44c: qq = 8'h2b; // 0x44c
	13'h44d: qq = 8'ha2; // 0x44d
	13'h44e: qq = 8'h2c; // 0x44e
	13'h44f: qq = 8'had; // 0x44f
	13'h450: qq = 8'h3c; // 0x450
	13'h451: qq = 8'hcb; // 0x451
	13'h452: qq = 8'h3c; // 0x452
	13'h453: qq = 8'he3; // 0x453
	13'h454: qq = 8'h3c; // 0x454
	13'h455: qq = 8'hfe; // 0x455
	13'h456: qq = 8'h3c; // 0x456
	13'h457: qq = 8'h19; // 0x457
	13'h458: qq = 8'h3d; // 0x458
	13'h459: qq = 8'h34; // 0x459
	13'h45a: qq = 8'h3d; // 0x45a
	13'h45b: qq = 8'h4f; // 0x45b
	13'h45c: qq = 8'h3d; // 0x45c
	13'h45d: qq = 8'h5d; // 0x45d
	13'h45e: qq = 8'h3d; // 0x45e
	13'h45f: qq = 8'h7d; // 0x45f
	13'h460: qq = 8'h3d; // 0x460
	13'h461: qq = 8'h9b; // 0x461
	13'h462: qq = 8'h3d; // 0x462
	13'h463: qq = 8'hbc; // 0x463
	13'h464: qq = 8'h3d; // 0x464
	13'h465: qq = 8'hdb; // 0x465
	13'h466: qq = 8'h3d; // 0x466
	13'h467: qq = 8'hf2; // 0x467
	13'h468: qq = 8'h3d; // 0x468
	13'h469: qq = 8'hf6; // 0x469
	13'h46a: qq = 8'h3d; // 0x46a
	13'h46b: qq = 8'hfd; // 0x46b
	13'h46c: qq = 8'h3d; // 0x46c
	13'h46d: qq = 8'h04; // 0x46d
	13'h46e: qq = 8'h3e; // 0x46e
	13'h46f: qq = 8'h0f; // 0x46f
	13'h470: qq = 8'h3e; // 0x470
	13'h471: qq = 8'ha0; // 0x471
	13'h472: qq = 8'h04; // 0x472
	13'h473: qq = 8'h40; // 0x473
	13'h474: qq = 8'h04; // 0x474
	13'h475: qq = 8'h20; // 0x475
	13'h476: qq = 8'h04; // 0x476
	13'h477: qq = 8'h60; // 0x477
	13'h478: qq = 8'h07; // 0x478
	13'h479: qq = 8'h60; // 0x479
	13'h47a: qq = 8'h07; // 0x47a
	13'h47b: qq = 8'h60; // 0x47b
	13'h47c: qq = 8'h07; // 0x47c
	13'h47d: qq = 8'h60; // 0x47d
	13'h47e: qq = 8'h07; // 0x47e
	13'h47f: qq = 8'he0; // 0x47f
	13'h480: qq = 8'h04; // 0x480
	13'h481: qq = 8'ha0; // 0x481
	13'h482: qq = 8'h04; // 0x482
	13'h483: qq = 8'h60; // 0x483
	13'h484: qq = 8'h07; // 0x484
	13'h485: qq = 8'he0; // 0x485
	13'h486: qq = 8'h04; // 0x486
	13'h487: qq = 8'h00; // 0x487
	13'h488: qq = 8'h04; // 0x488
	13'h489: qq = 8'h75; // 0x489
	13'h48a: qq = 8'h07; // 0x48a
	13'h48b: qq = 8'h75; // 0x48b
	13'h48c: qq = 8'h07; // 0x48c
	13'h48d: qq = 8'h75; // 0x48d
	13'h48e: qq = 8'h07; // 0x48e
	13'h48f: qq = 8'h6b; // 0x48f
	13'h490: qq = 8'h04; // 0x490
	13'h491: qq = 8'h2e; // 0x491
	13'h492: qq = 8'h04; // 0x492
	13'h493: qq = 8'h40; // 0x493
	13'h494: qq = 8'h04; // 0x494
	13'h495: qq = 8'h60; // 0x495
	13'h496: qq = 8'h04; // 0x496
	13'h497: qq = 8'h80; // 0x497
	13'h498: qq = 8'h04; // 0x498
	13'h499: qq = 8'ha0; // 0x499
	13'h49a: qq = 8'h04; // 0x49a
	13'h49b: qq = 8'hc0; // 0x49b
	13'h49c: qq = 8'h04; // 0x49c
	13'h49d: qq = 8'he0; // 0x49d
	13'h49e: qq = 8'h04; // 0x49e
	13'h49f: qq = 8'h00; // 0x49f
	13'h4a0: qq = 8'h05; // 0x4a0
	13'h4a1: qq = 8'h0c; // 0x4a1
	13'h4a2: qq = 8'h08; // 0x4a2
	13'h4a3: qq = 8'h06; // 0x4a3
	13'h4a4: qq = 8'h05; // 0x4a4
	13'h4a5: qq = 8'h26; // 0x4a5
	13'h4a6: qq = 8'h38; // 0x4a6
	13'h4a7: qq = 8'h4b; // 0x4a7
	13'h4a8: qq = 8'h5e; // 0x4a8
	13'h4a9: qq = 8'ha0; // 0x4a9
	13'h4aa: qq = 8'h90; // 0x4aa
	13'h4ab: qq = 8'h80; // 0x4ab
	13'h4ac: qq = 8'h70; // 0x4ac
	13'h4ad: qq = 8'h20; // 0x4ad
	13'h4ae: qq = 8'h20; // 0x4ae
	13'h4af: qq = 8'h20; // 0x4af
	13'h4b0: qq = 8'h20; // 0x4b0
	13'h4b1: qq = 8'h20; // 0x4b1
	13'h4b2: qq = 8'h20; // 0x4b2
	13'h4b3: qq = 8'h20; // 0x4b3
	13'h4b4: qq = 8'h59; // 0x4b4
	13'h4b5: qq = 8'h4f; // 0x4b5
	13'h4b6: qq = 8'h55; // 0x4b6
	13'h4b7: qq = 8'h52; // 0x4b7
	13'h4b8: qq = 8'h20; // 0x4b8
	13'h4b9: qq = 8'h43; // 0x4b9
	13'h4ba: qq = 8'h41; // 0x4ba
	13'h4bb: qq = 8'h52; // 0x4bb
	13'h4bc: qq = 8'h20; // 0x4bc
	13'h4bd: qq = 8'h49; // 0x4bd
	13'h4be: qq = 8'h53; // 0x4be
	13'h4bf: qq = 8'h20; // 0x4bf
	13'h4c0: qq = 8'hd7; // 0x4c0
	13'h4c1: qq = 8'hc8; // 0x4c1
	13'h4c2: qq = 8'hc9; // 0x4c2
	13'h4c3: qq = 8'hd4; // 0x4c3
	13'h4c4: qq = 8'hc5; // 0x4c4
	13'h4c5: qq = 8'h20; // 0x4c5
	13'h4c6: qq = 8'h20; // 0x4c6
	13'h4c7: qq = 8'h20; // 0x4c7
	13'h4c8: qq = 8'h20; // 0x4c8
	13'h4c9: qq = 8'h20; // 0x4c9
	13'h4ca: qq = 8'h00; // 0x4ca
	13'h4cb: qq = 8'h20; // 0x4cb
	13'h4cc: qq = 8'h20; // 0x4cc
	13'h4cd: qq = 8'h20; // 0x4cd
	13'h4ce: qq = 8'h20; // 0x4ce
	13'h4cf: qq = 8'h20; // 0x4cf
	13'h4d0: qq = 8'h20; // 0x4d0
	13'h4d1: qq = 8'h20; // 0x4d1
	13'h4d2: qq = 8'h20; // 0x4d2
	13'h4d3: qq = 8'h20; // 0x4d3
	13'h4d4: qq = 8'h20; // 0x4d4
	13'h4d5: qq = 8'h45; // 0x4d5
	13'h4d6: qq = 8'h58; // 0x4d6
	13'h4d7: qq = 8'h54; // 0x4d7
	13'h4d8: qq = 8'h45; // 0x4d8
	13'h4d9: qq = 8'h4e; // 0x4d9
	13'h4da: qq = 8'h44; // 0x4da
	13'h4db: qq = 8'h45; // 0x4db
	13'h4dc: qq = 8'h44; // 0x4dc
	13'h4dd: qq = 8'h20; // 0x4dd
	13'h4de: qq = 8'h50; // 0x4de
	13'h4df: qq = 8'h4c; // 0x4df
	13'h4e0: qq = 8'h41; // 0x4e0
	13'h4e1: qq = 8'h59; // 0x4e1
	13'h4e2: qq = 8'h00; // 0x4e2
	13'h4e3: qq = 8'h20; // 0x4e3
	13'h4e4: qq = 8'h20; // 0x4e4
	13'h4e5: qq = 8'h53; // 0x4e5
	13'h4e6: qq = 8'h43; // 0x4e6
	13'h4e7: qq = 8'h4f; // 0x4e7
	13'h4e8: qq = 8'h52; // 0x4e8
	13'h4e9: qq = 8'h45; // 0x4e9
	13'h4ea: qq = 8'h20; // 0x4ea
	13'h4eb: qq = 8'h20; // 0x4eb
	13'h4ec: qq = 8'h20; // 0x4ec
	13'h4ed: qq = 8'h20; // 0x4ed
	13'h4ee: qq = 8'h20; // 0x4ee
	13'h4ef: qq = 8'h20; // 0x4ef
	13'h4f0: qq = 8'h20; // 0x4f0
	13'h4f1: qq = 8'h20; // 0x4f1
	13'h4f2: qq = 8'h20; // 0x4f2
	13'h4f3: qq = 8'h20; // 0x4f3
	13'h4f4: qq = 8'h20; // 0x4f4
	13'h4f5: qq = 8'h20; // 0x4f5
	13'h4f6: qq = 8'h20; // 0x4f6
	13'h4f7: qq = 8'h20; // 0x4f7
	13'h4f8: qq = 8'h54; // 0x4f8
	13'h4f9: qq = 8'h49; // 0x4f9
	13'h4fa: qq = 8'h4d; // 0x4fa
	13'h4fb: qq = 8'h45; // 0x4fb
	13'h4fc: qq = 8'h20; // 0x4fc
	13'h4fd: qq = 8'h00; // 0x4fd
	13'h4fe: qq = 8'h20; // 0x4fe
	13'h4ff: qq = 8'h20; // 0x4ff
	13'h500: qq = 8'h20; // 0x500
	13'h501: qq = 8'h20; // 0x501
	13'h502: qq = 8'h20; // 0x502
	13'h503: qq = 8'h20; // 0x503
	13'h504: qq = 8'h20; // 0x504
	13'h505: qq = 8'h20; // 0x505
	13'h506: qq = 8'h31; // 0x506
	13'h507: qq = 8'h20; // 0x507
	13'h508: qq = 8'h43; // 0x508
	13'h509: qq = 8'h4f; // 0x509
	13'h50a: qq = 8'h49; // 0x50a
	13'h50b: qq = 8'h4e; // 0x50b
	13'h50c: qq = 8'h20; // 0x50c
	13'h50d: qq = 8'h50; // 0x50d
	13'h50e: qq = 8'h45; // 0x50e
	13'h50f: qq = 8'h52; // 0x50f
	13'h510: qq = 8'h20; // 0x510
	13'h511: qq = 8'h47; // 0x511
	13'h512: qq = 8'h41; // 0x512
	13'h513: qq = 8'h4d; // 0x513
	13'h514: qq = 8'h45; // 0x514
	13'h515: qq = 8'h20; // 0x515
	13'h516: qq = 8'h20; // 0x516
	13'h517: qq = 8'h20; // 0x517
	13'h518: qq = 8'h00; // 0x518
	13'h519: qq = 8'h20; // 0x519
	13'h51a: qq = 8'h20; // 0x51a
	13'h51b: qq = 8'h20; // 0x51b
	13'h51c: qq = 8'h20; // 0x51c
	13'h51d: qq = 8'h20; // 0x51d
	13'h51e: qq = 8'h20; // 0x51e
	13'h51f: qq = 8'h20; // 0x51f
	13'h520: qq = 8'h32; // 0x520
	13'h521: qq = 8'h20; // 0x521
	13'h522: qq = 8'h43; // 0x522
	13'h523: qq = 8'h4f; // 0x523
	13'h524: qq = 8'h49; // 0x524
	13'h525: qq = 8'h4e; // 0x525
	13'h526: qq = 8'h53; // 0x526
	13'h527: qq = 8'h20; // 0x527
	13'h528: qq = 8'h50; // 0x528
	13'h529: qq = 8'h45; // 0x529
	13'h52a: qq = 8'h52; // 0x52a
	13'h52b: qq = 8'h20; // 0x52b
	13'h52c: qq = 8'h47; // 0x52c
	13'h52d: qq = 8'h41; // 0x52d
	13'h52e: qq = 8'h4d; // 0x52e
	13'h52f: qq = 8'h45; // 0x52f
	13'h530: qq = 8'h20; // 0x530
	13'h531: qq = 8'h20; // 0x531
	13'h532: qq = 8'h20; // 0x532
	13'h533: qq = 8'h00; // 0x533
	13'h534: qq = 8'h20; // 0x534
	13'h535: qq = 8'h20; // 0x535
	13'h536: qq = 8'h20; // 0x536
	13'h537: qq = 8'h20; // 0x537
	13'h538: qq = 8'h20; // 0x538
	13'h539: qq = 8'h20; // 0x539
	13'h53a: qq = 8'h20; // 0x53a
	13'h53b: qq = 8'h20; // 0x53b
	13'h53c: qq = 8'h32; // 0x53c
	13'h53d: qq = 8'h20; // 0x53d
	13'h53e: qq = 8'h47; // 0x53e
	13'h53f: qq = 8'h41; // 0x53f
	13'h540: qq = 8'h4d; // 0x540
	13'h541: qq = 8'h45; // 0x541
	13'h542: qq = 8'h53; // 0x542
	13'h543: qq = 8'h20; // 0x543
	13'h544: qq = 8'h50; // 0x544
	13'h545: qq = 8'h45; // 0x545
	13'h546: qq = 8'h52; // 0x546
	13'h547: qq = 8'h20; // 0x547
	13'h548: qq = 8'h43; // 0x548
	13'h549: qq = 8'h4f; // 0x549
	13'h54a: qq = 8'h49; // 0x54a
	13'h54b: qq = 8'h4e; // 0x54b
	13'h54c: qq = 8'h20; // 0x54c
	13'h54d: qq = 8'h20; // 0x54d
	13'h54e: qq = 8'h00; // 0x54e
	13'h54f: qq = 8'h20; // 0x54f
	13'h550: qq = 8'h20; // 0x550
	13'h551: qq = 8'h20; // 0x551
	13'h552: qq = 8'h20; // 0x552
	13'h553: qq = 8'h20; // 0x553
	13'h554: qq = 8'h20; // 0x554
	13'h555: qq = 8'h20; // 0x555
	13'h556: qq = 8'h52; // 0x556
	13'h557: qq = 8'h41; // 0x557
	13'h558: qq = 8'h54; // 0x558
	13'h559: qq = 8'h49; // 0x559
	13'h55a: qq = 8'h4e; // 0x55a
	13'h55b: qq = 8'h47; // 0x55b
	13'h55c: qq = 8'h00; // 0x55c
	13'h55d: qq = 8'h20; // 0x55d
	13'h55e: qq = 8'h42; // 0x55e
	13'h55f: qq = 8'h4c; // 0x55f
	13'h560: qq = 8'h41; // 0x560
	13'h561: qq = 8'h43; // 0x561
	13'h562: qq = 8'h4b; // 0x562
	13'h563: qq = 8'h20; // 0x563
	13'h564: qq = 8'h43; // 0x564
	13'h565: qq = 8'h41; // 0x565
	13'h566: qq = 8'h52; // 0x566
	13'h567: qq = 8'h53; // 0x567
	13'h568: qq = 8'h20; // 0x568
	13'h569: qq = 8'h44; // 0x569
	13'h56a: qq = 8'h52; // 0x56a
	13'h56b: qq = 8'h49; // 0x56b
	13'h56c: qq = 8'h56; // 0x56c
	13'h56d: qq = 8'h45; // 0x56d
	13'h56e: qq = 8'h20; // 0x56e
	13'h56f: qq = 8'h41; // 0x56f
	13'h570: qq = 8'h55; // 0x570
	13'h571: qq = 8'h54; // 0x571
	13'h572: qq = 8'h4f; // 0x572
	13'h573: qq = 8'h4d; // 0x573
	13'h574: qq = 8'h41; // 0x574
	13'h575: qq = 8'h54; // 0x575
	13'h576: qq = 8'h49; // 0x576
	13'h577: qq = 8'h43; // 0x577
	13'h578: qq = 8'h41; // 0x578
	13'h579: qq = 8'h4c; // 0x579
	13'h57a: qq = 8'h4c; // 0x57a
	13'h57b: qq = 8'h59; // 0x57b
	13'h57c: qq = 8'h00; // 0x57c
	13'h57d: qq = 8'h20; // 0x57d
	13'h57e: qq = 8'h20; // 0x57e
	13'h57f: qq = 8'h54; // 0x57f
	13'h580: qq = 8'h52; // 0x580
	13'h581: qq = 8'h41; // 0x581
	13'h582: qq = 8'h43; // 0x582
	13'h583: qq = 8'h4b; // 0x583
	13'h584: qq = 8'h53; // 0x584
	13'h585: qq = 8'h20; // 0x585
	13'h586: qq = 8'h43; // 0x586
	13'h587: qq = 8'h48; // 0x587
	13'h588: qq = 8'h41; // 0x588
	13'h589: qq = 8'h4e; // 0x589
	13'h58a: qq = 8'h47; // 0x58a
	13'h58b: qq = 8'h45; // 0x58b
	13'h58c: qq = 8'h20; // 0x58c
	13'h58d: qq = 8'h41; // 0x58d
	13'h58e: qq = 8'h55; // 0x58e
	13'h58f: qq = 8'h54; // 0x58f
	13'h590: qq = 8'h4f; // 0x590
	13'h591: qq = 8'h4d; // 0x591
	13'h592: qq = 8'h41; // 0x592
	13'h593: qq = 8'h54; // 0x593
	13'h594: qq = 8'h49; // 0x594
	13'h595: qq = 8'h43; // 0x595
	13'h596: qq = 8'h41; // 0x596
	13'h597: qq = 8'h4c; // 0x597
	13'h598: qq = 8'h4c; // 0x598
	13'h599: qq = 8'h59; // 0x599
	13'h59a: qq = 8'h00; // 0x59a
	13'h59b: qq = 8'h20; // 0x59b
	13'h59c: qq = 8'h20; // 0x59c
	13'h59d: qq = 8'h45; // 0x59d
	13'h59e: qq = 8'h58; // 0x59e
	13'h59f: qq = 8'h54; // 0x59f
	13'h5a0: qq = 8'h45; // 0x5a0
	13'h5a1: qq = 8'h4e; // 0x5a1
	13'h5a2: qq = 8'h44; // 0x5a2
	13'h5a3: qq = 8'h45; // 0x5a3
	13'h5a4: qq = 8'h44; // 0x5a4
	13'h5a5: qq = 8'h20; // 0x5a5
	13'h5a6: qq = 8'h50; // 0x5a6
	13'h5a7: qq = 8'h4c; // 0x5a7
	13'h5a8: qq = 8'h41; // 0x5a8
	13'h5a9: qq = 8'h59; // 0x5a9
	13'h5aa: qq = 8'h20; // 0x5aa
	13'h5ab: qq = 8'h46; // 0x5ab
	13'h5ac: qq = 8'h4f; // 0x5ac
	13'h5ad: qq = 8'h52; // 0x5ad
	13'h5ae: qq = 8'h20; // 0x5ae
	13'h5af: qq = 8'h20; // 0x5af
	13'h5b0: qq = 8'h20; // 0x5b0
	13'h5b1: qq = 8'h30; // 0x5b1
	13'h5b2: qq = 8'h20; // 0x5b2
	13'h5b3: qq = 8'h50; // 0x5b3
	13'h5b4: qq = 8'h4f; // 0x5b4
	13'h5b5: qq = 8'h49; // 0x5b5
	13'h5b6: qq = 8'h4e; // 0x5b6
	13'h5b7: qq = 8'h54; // 0x5b7
	13'h5b8: qq = 8'h53; // 0x5b8
	13'h5b9: qq = 8'h20; // 0x5b9
	13'h5ba: qq = 8'h20; // 0x5ba
	13'h5bb: qq = 8'h00; // 0x5bb
	13'h5bc: qq = 8'h20; // 0x5bc
	13'h5bd: qq = 8'h20; // 0x5bd
	13'h5be: qq = 8'h20; // 0x5be
	13'h5bf: qq = 8'h20; // 0x5bf
	13'h5c0: qq = 8'h20; // 0x5c0
	13'h5c1: qq = 8'h20; // 0x5c1
	13'h5c2: qq = 8'h20; // 0x5c2
	13'h5c3: qq = 8'h50; // 0x5c3
	13'h5c4: qq = 8'h55; // 0x5c4
	13'h5c5: qq = 8'h53; // 0x5c5
	13'h5c6: qq = 8'h48; // 0x5c6
	13'h5c7: qq = 8'h20; // 0x5c7
	13'h5c8: qq = 8'h53; // 0x5c8
	13'h5c9: qq = 8'h54; // 0x5c9
	13'h5ca: qq = 8'h41; // 0x5ca
	13'h5cb: qq = 8'h52; // 0x5cb
	13'h5cc: qq = 8'h54; // 0x5cc
	13'h5cd: qq = 8'h20; // 0x5cd
	13'h5ce: qq = 8'h42; // 0x5ce
	13'h5cf: qq = 8'h55; // 0x5cf
	13'h5d0: qq = 8'h54; // 0x5d0
	13'h5d1: qq = 8'h54; // 0x5d1
	13'h5d2: qq = 8'h4f; // 0x5d2
	13'h5d3: qq = 8'h4e; // 0x5d3
	13'h5d4: qq = 8'h20; // 0x5d4
	13'h5d5: qq = 8'h20; // 0x5d5
	13'h5d6: qq = 8'h20; // 0x5d6
	13'h5d7: qq = 8'h20; // 0x5d7
	13'h5d8: qq = 8'h20; // 0x5d8
	13'h5d9: qq = 8'h20; // 0x5d9
	13'h5da: qq = 8'h00; // 0x5da
	13'h5db: qq = 8'h20; // 0x5db
	13'h5dc: qq = 8'h20; // 0x5dc
	13'h5dd: qq = 8'h20; // 0x5dd
	13'h5de: qq = 8'h20; // 0x5de
	13'h5df: qq = 8'h20; // 0x5df
	13'h5e0: qq = 8'h20; // 0x5e0
	13'h5e1: qq = 8'h20; // 0x5e1
	13'h5e2: qq = 8'h20; // 0x5e2
	13'h5e3: qq = 8'h20; // 0x5e3
	13'h5e4: qq = 8'h20; // 0x5e4
	13'h5e5: qq = 8'h20; // 0x5e5
	13'h5e6: qq = 8'h20; // 0x5e6
	13'h5e7: qq = 8'h47; // 0x5e7
	13'h5e8: qq = 8'h41; // 0x5e8
	13'h5e9: qq = 8'h4d; // 0x5e9
	13'h5ea: qq = 8'h45; // 0x5ea
	13'h5eb: qq = 8'h20; // 0x5eb
	13'h5ec: qq = 8'h20; // 0x5ec
	13'h5ed: qq = 8'h4f; // 0x5ed
	13'h5ee: qq = 8'h56; // 0x5ee
	13'h5ef: qq = 8'h45; // 0x5ef
	13'h5f0: qq = 8'h52; // 0x5f0
	13'h5f1: qq = 8'h00; // 0x5f1
	13'h5f2: qq = 8'h50; // 0x5f2
	13'h5f3: qq = 8'h52; // 0x5f3
	13'h5f4: qq = 8'h4f; // 0x5f4
	13'h5f5: qq = 8'h00; // 0x5f5
	13'h5f6: qq = 8'h52; // 0x5f6
	13'h5f7: qq = 8'h4f; // 0x5f7
	13'h5f8: qq = 8'h4f; // 0x5f8
	13'h5f9: qq = 8'h4b; // 0x5f9
	13'h5fa: qq = 8'h49; // 0x5fa
	13'h5fb: qq = 8'h45; // 0x5fb
	13'h5fc: qq = 8'h00; // 0x5fc
	13'h5fd: qq = 8'h47; // 0x5fd
	13'h5fe: qq = 8'h52; // 0x5fe
	13'h5ff: qq = 8'h41; // 0x5ff
	13'h600: qq = 8'h4e; // 0x600
	13'h601: qq = 8'h4e; // 0x601
	13'h602: qq = 8'h59; // 0x602
	13'h603: qq = 8'h00; // 0x603
	13'h604: qq = 8'h4b; // 0x604
	13'h605: qq = 8'h45; // 0x605
	13'h606: qq = 8'h45; // 0x606
	13'h607: qq = 8'h20; // 0x607
	13'h608: qq = 8'h20; // 0x608
	13'h609: qq = 8'h47; // 0x609
	13'h60a: qq = 8'h41; // 0x60a
	13'h60b: qq = 8'h4d; // 0x60b
	13'h60c: qq = 8'h45; // 0x60c
	13'h60d: qq = 8'h53; // 0x60d
	13'h60e: qq = 8'h00; // 0x60e
	13'h60f: qq = 8'h48; // 0x60f
	13'h610: qq = 8'h49; // 0x610
	13'h611: qq = 8'h47; // 0x611
	13'h612: qq = 8'h48; // 0x612
	13'h613: qq = 8'h20; // 0x613
	13'h614: qq = 8'h53; // 0x614
	13'h615: qq = 8'h43; // 0x615
	13'h616: qq = 8'h4f; // 0x616
	13'h617: qq = 8'h52; // 0x617
	13'h618: qq = 8'h45; // 0x618
	13'h619: qq = 8'h20; // 0x619
	13'h61a: qq = 8'h20; // 0x61a
	13'h61b: qq = 8'h20; // 0x61b
	13'h61c: qq = 8'h20; // 0x61c
	13'h61d: qq = 8'h20; // 0x61d
	13'h61e: qq = 8'h00; // 0x61e
	13'h61f: qq = 8'h00; // 0x61f
	13'h620: qq = 8'h00; // 0x620
	13'h621: qq = 8'h00; // 0x621
	13'h622: qq = 8'h00; // 0x622
	13'h623: qq = 8'h00; // 0x623
	13'h624: qq = 8'h00; // 0x624
	13'h625: qq = 8'h00; // 0x625
	13'h626: qq = 8'h00; // 0x626
	13'h627: qq = 8'h00; // 0x627
	13'h628: qq = 8'h00; // 0x628
	13'h629: qq = 8'h00; // 0x629
	13'h62a: qq = 8'h00; // 0x62a
	13'h62b: qq = 8'h00; // 0x62b
	13'h62c: qq = 8'h00; // 0x62c
	13'h62d: qq = 8'h00; // 0x62d
	13'h62e: qq = 8'h00; // 0x62e
	13'h62f: qq = 8'h00; // 0x62f
	13'h630: qq = 8'h00; // 0x630
	13'h631: qq = 8'h00; // 0x631
	13'h632: qq = 8'h00; // 0x632
	13'h633: qq = 8'h00; // 0x633
	13'h634: qq = 8'h00; // 0x634
	13'h635: qq = 8'h00; // 0x635
	13'h636: qq = 8'h00; // 0x636
	13'h637: qq = 8'h00; // 0x637
	13'h638: qq = 8'h00; // 0x638
	13'h639: qq = 8'h00; // 0x639
	13'h63a: qq = 8'h00; // 0x63a
	13'h63b: qq = 8'h00; // 0x63b
	13'h63c: qq = 8'h00; // 0x63c
	13'h63d: qq = 8'h00; // 0x63d
	13'h63e: qq = 8'h00; // 0x63e
	13'h63f: qq = 8'h00; // 0x63f
	13'h640: qq = 8'h00; // 0x640
	13'h641: qq = 8'h00; // 0x641
	13'h642: qq = 8'h00; // 0x642
	13'h643: qq = 8'h00; // 0x643
	13'h644: qq = 8'h00; // 0x644
	13'h645: qq = 8'h00; // 0x645
	13'h646: qq = 8'h00; // 0x646
	13'h647: qq = 8'h00; // 0x647
	13'h648: qq = 8'h00; // 0x648
	13'h649: qq = 8'h00; // 0x649
	13'h64a: qq = 8'h00; // 0x64a
	13'h64b: qq = 8'h00; // 0x64b
	13'h64c: qq = 8'h00; // 0x64c
	13'h64d: qq = 8'h00; // 0x64d
	13'h64e: qq = 8'h00; // 0x64e
	13'h64f: qq = 8'h00; // 0x64f
	13'h650: qq = 8'h00; // 0x650
	13'h651: qq = 8'h00; // 0x651
	13'h652: qq = 8'h00; // 0x652
	13'h653: qq = 8'h00; // 0x653
	13'h654: qq = 8'h00; // 0x654
	13'h655: qq = 8'h00; // 0x655
	13'h656: qq = 8'h00; // 0x656
	13'h657: qq = 8'h00; // 0x657
	13'h658: qq = 8'h00; // 0x658
	13'h659: qq = 8'h00; // 0x659
	13'h65a: qq = 8'h00; // 0x65a
	13'h65b: qq = 8'h00; // 0x65b
	13'h65c: qq = 8'h00; // 0x65c
	13'h65d: qq = 8'h00; // 0x65d
	13'h65e: qq = 8'h00; // 0x65e
	13'h65f: qq = 8'h00; // 0x65f
	13'h660: qq = 8'h00; // 0x660
	13'h661: qq = 8'h00; // 0x661
	13'h662: qq = 8'h00; // 0x662
	13'h663: qq = 8'h00; // 0x663
	13'h664: qq = 8'h00; // 0x664
	13'h665: qq = 8'h00; // 0x665
	13'h666: qq = 8'h00; // 0x666
	13'h667: qq = 8'h00; // 0x667
	13'h668: qq = 8'h00; // 0x668
	13'h669: qq = 8'h00; // 0x669
	13'h66a: qq = 8'h00; // 0x66a
	13'h66b: qq = 8'h00; // 0x66b
	13'h66c: qq = 8'h00; // 0x66c
	13'h66d: qq = 8'h00; // 0x66d
	13'h66e: qq = 8'h00; // 0x66e
	13'h66f: qq = 8'h00; // 0x66f
	13'h670: qq = 8'h00; // 0x670
	13'h671: qq = 8'h00; // 0x671
	13'h672: qq = 8'h00; // 0x672
	13'h673: qq = 8'h00; // 0x673
	13'h674: qq = 8'h00; // 0x674
	13'h675: qq = 8'h00; // 0x675
	13'h676: qq = 8'h00; // 0x676
	13'h677: qq = 8'h00; // 0x677
	13'h678: qq = 8'h00; // 0x678
	13'h679: qq = 8'h00; // 0x679
	13'h67a: qq = 8'h00; // 0x67a
	13'h67b: qq = 8'h00; // 0x67b
	13'h67c: qq = 8'h00; // 0x67c
	13'h67d: qq = 8'h00; // 0x67d
	13'h67e: qq = 8'h00; // 0x67e
	13'h67f: qq = 8'h00; // 0x67f
	13'h680: qq = 8'h00; // 0x680
	13'h681: qq = 8'h00; // 0x681
	13'h682: qq = 8'h00; // 0x682
	13'h683: qq = 8'h00; // 0x683
	13'h684: qq = 8'h00; // 0x684
	13'h685: qq = 8'h00; // 0x685
	13'h686: qq = 8'h00; // 0x686
	13'h687: qq = 8'h00; // 0x687
	13'h688: qq = 8'h00; // 0x688
	13'h689: qq = 8'h00; // 0x689
	13'h68a: qq = 8'h00; // 0x68a
	13'h68b: qq = 8'h00; // 0x68b
	13'h68c: qq = 8'h00; // 0x68c
	13'h68d: qq = 8'h00; // 0x68d
	13'h68e: qq = 8'h00; // 0x68e
	13'h68f: qq = 8'h00; // 0x68f
	13'h690: qq = 8'h00; // 0x690
	13'h691: qq = 8'h00; // 0x691
	13'h692: qq = 8'h00; // 0x692
	13'h693: qq = 8'h00; // 0x693
	13'h694: qq = 8'h00; // 0x694
	13'h695: qq = 8'h00; // 0x695
	13'h696: qq = 8'h00; // 0x696
	13'h697: qq = 8'h00; // 0x697
	13'h698: qq = 8'h00; // 0x698
	13'h699: qq = 8'h00; // 0x699
	13'h69a: qq = 8'h00; // 0x69a
	13'h69b: qq = 8'h00; // 0x69b
	13'h69c: qq = 8'h00; // 0x69c
	13'h69d: qq = 8'h00; // 0x69d
	13'h69e: qq = 8'h00; // 0x69e
	13'h69f: qq = 8'h00; // 0x69f
	13'h6a0: qq = 8'h00; // 0x6a0
	13'h6a1: qq = 8'h00; // 0x6a1
	13'h6a2: qq = 8'h00; // 0x6a2
	13'h6a3: qq = 8'h00; // 0x6a3
	13'h6a4: qq = 8'h00; // 0x6a4
	13'h6a5: qq = 8'h00; // 0x6a5
	13'h6a6: qq = 8'h00; // 0x6a6
	13'h6a7: qq = 8'h00; // 0x6a7
	13'h6a8: qq = 8'h00; // 0x6a8
	13'h6a9: qq = 8'h00; // 0x6a9
	13'h6aa: qq = 8'h00; // 0x6aa
	13'h6ab: qq = 8'h00; // 0x6ab
	13'h6ac: qq = 8'h00; // 0x6ac
	13'h6ad: qq = 8'h00; // 0x6ad
	13'h6ae: qq = 8'h00; // 0x6ae
	13'h6af: qq = 8'h00; // 0x6af
	13'h6b0: qq = 8'h00; // 0x6b0
	13'h6b1: qq = 8'h00; // 0x6b1
	13'h6b2: qq = 8'h00; // 0x6b2
	13'h6b3: qq = 8'h00; // 0x6b3
	13'h6b4: qq = 8'h00; // 0x6b4
	13'h6b5: qq = 8'h00; // 0x6b5
	13'h6b6: qq = 8'h00; // 0x6b6
	13'h6b7: qq = 8'h00; // 0x6b7
	13'h6b8: qq = 8'h00; // 0x6b8
	13'h6b9: qq = 8'h00; // 0x6b9
	13'h6ba: qq = 8'h00; // 0x6ba
	13'h6bb: qq = 8'h00; // 0x6bb
	13'h6bc: qq = 8'h00; // 0x6bc
	13'h6bd: qq = 8'h00; // 0x6bd
	13'h6be: qq = 8'h00; // 0x6be
	13'h6bf: qq = 8'h00; // 0x6bf
	13'h6c0: qq = 8'h00; // 0x6c0
	13'h6c1: qq = 8'h00; // 0x6c1
	13'h6c2: qq = 8'h00; // 0x6c2
	13'h6c3: qq = 8'h00; // 0x6c3
	13'h6c4: qq = 8'h00; // 0x6c4
	13'h6c5: qq = 8'h00; // 0x6c5
	13'h6c6: qq = 8'h00; // 0x6c6
	13'h6c7: qq = 8'h00; // 0x6c7
	13'h6c8: qq = 8'h00; // 0x6c8
	13'h6c9: qq = 8'h00; // 0x6c9
	13'h6ca: qq = 8'h00; // 0x6ca
	13'h6cb: qq = 8'h00; // 0x6cb
	13'h6cc: qq = 8'h00; // 0x6cc
	13'h6cd: qq = 8'h00; // 0x6cd
	13'h6ce: qq = 8'h00; // 0x6ce
	13'h6cf: qq = 8'h00; // 0x6cf
	13'h6d0: qq = 8'h00; // 0x6d0
	13'h6d1: qq = 8'h00; // 0x6d1
	13'h6d2: qq = 8'h00; // 0x6d2
	13'h6d3: qq = 8'h00; // 0x6d3
	13'h6d4: qq = 8'h00; // 0x6d4
	13'h6d5: qq = 8'h00; // 0x6d5
	13'h6d6: qq = 8'h00; // 0x6d6
	13'h6d7: qq = 8'h00; // 0x6d7
	13'h6d8: qq = 8'h00; // 0x6d8
	13'h6d9: qq = 8'h00; // 0x6d9
	13'h6da: qq = 8'h00; // 0x6da
	13'h6db: qq = 8'h00; // 0x6db
	13'h6dc: qq = 8'h00; // 0x6dc
	13'h6dd: qq = 8'h00; // 0x6dd
	13'h6de: qq = 8'h00; // 0x6de
	13'h6df: qq = 8'h00; // 0x6df
	13'h6e0: qq = 8'h00; // 0x6e0
	13'h6e1: qq = 8'h00; // 0x6e1
	13'h6e2: qq = 8'h00; // 0x6e2
	13'h6e3: qq = 8'h00; // 0x6e3
	13'h6e4: qq = 8'h00; // 0x6e4
	13'h6e5: qq = 8'h00; // 0x6e5
	13'h6e6: qq = 8'h00; // 0x6e6
	13'h6e7: qq = 8'h00; // 0x6e7
	13'h6e8: qq = 8'h00; // 0x6e8
	13'h6e9: qq = 8'h00; // 0x6e9
	13'h6ea: qq = 8'h00; // 0x6ea
	13'h6eb: qq = 8'h00; // 0x6eb
	13'h6ec: qq = 8'h00; // 0x6ec
	13'h6ed: qq = 8'h00; // 0x6ed
	13'h6ee: qq = 8'h00; // 0x6ee
	13'h6ef: qq = 8'h00; // 0x6ef
	13'h6f0: qq = 8'h00; // 0x6f0
	13'h6f1: qq = 8'h00; // 0x6f1
	13'h6f2: qq = 8'h00; // 0x6f2
	13'h6f3: qq = 8'h00; // 0x6f3
	13'h6f4: qq = 8'h00; // 0x6f4
	13'h6f5: qq = 8'h00; // 0x6f5
	13'h6f6: qq = 8'h00; // 0x6f6
	13'h6f7: qq = 8'h00; // 0x6f7
	13'h6f8: qq = 8'h00; // 0x6f8
	13'h6f9: qq = 8'h00; // 0x6f9
	13'h6fa: qq = 8'h00; // 0x6fa
	13'h6fb: qq = 8'h00; // 0x6fb
	13'h6fc: qq = 8'h00; // 0x6fc
	13'h6fd: qq = 8'h00; // 0x6fd
	13'h6fe: qq = 8'h00; // 0x6fe
	13'h6ff: qq = 8'h00; // 0x6ff
	13'h700: qq = 8'h00; // 0x700
	13'h701: qq = 8'h00; // 0x701
	13'h702: qq = 8'h00; // 0x702
	13'h703: qq = 8'h00; // 0x703
	13'h704: qq = 8'h00; // 0x704
	13'h705: qq = 8'h00; // 0x705
	13'h706: qq = 8'h00; // 0x706
	13'h707: qq = 8'h00; // 0x707
	13'h708: qq = 8'h00; // 0x708
	13'h709: qq = 8'h00; // 0x709
	13'h70a: qq = 8'h00; // 0x70a
	13'h70b: qq = 8'h00; // 0x70b
	13'h70c: qq = 8'h00; // 0x70c
	13'h70d: qq = 8'h00; // 0x70d
	13'h70e: qq = 8'h00; // 0x70e
	13'h70f: qq = 8'h00; // 0x70f
	13'h710: qq = 8'h00; // 0x710
	13'h711: qq = 8'h00; // 0x711
	13'h712: qq = 8'h00; // 0x712
	13'h713: qq = 8'h00; // 0x713
	13'h714: qq = 8'h00; // 0x714
	13'h715: qq = 8'h00; // 0x715
	13'h716: qq = 8'h00; // 0x716
	13'h717: qq = 8'h00; // 0x717
	13'h718: qq = 8'h00; // 0x718
	13'h719: qq = 8'h00; // 0x719
	13'h71a: qq = 8'h00; // 0x71a
	13'h71b: qq = 8'h00; // 0x71b
	13'h71c: qq = 8'h00; // 0x71c
	13'h71d: qq = 8'h00; // 0x71d
	13'h71e: qq = 8'h00; // 0x71e
	13'h71f: qq = 8'h00; // 0x71f
	13'h720: qq = 8'h00; // 0x720
	13'h721: qq = 8'h00; // 0x721
	13'h722: qq = 8'h00; // 0x722
	13'h723: qq = 8'h00; // 0x723
	13'h724: qq = 8'h00; // 0x724
	13'h725: qq = 8'h00; // 0x725
	13'h726: qq = 8'h00; // 0x726
	13'h727: qq = 8'h00; // 0x727
	13'h728: qq = 8'h00; // 0x728
	13'h729: qq = 8'h00; // 0x729
	13'h72a: qq = 8'h00; // 0x72a
	13'h72b: qq = 8'h00; // 0x72b
	13'h72c: qq = 8'h00; // 0x72c
	13'h72d: qq = 8'h00; // 0x72d
	13'h72e: qq = 8'h00; // 0x72e
	13'h72f: qq = 8'h00; // 0x72f
	13'h730: qq = 8'h00; // 0x730
	13'h731: qq = 8'h00; // 0x731
	13'h732: qq = 8'h00; // 0x732
	13'h733: qq = 8'h00; // 0x733
	13'h734: qq = 8'h00; // 0x734
	13'h735: qq = 8'h00; // 0x735
	13'h736: qq = 8'h00; // 0x736
	13'h737: qq = 8'h00; // 0x737
	13'h738: qq = 8'h00; // 0x738
	13'h739: qq = 8'h00; // 0x739
	13'h73a: qq = 8'h00; // 0x73a
	13'h73b: qq = 8'h00; // 0x73b
	13'h73c: qq = 8'h00; // 0x73c
	13'h73d: qq = 8'h00; // 0x73d
	13'h73e: qq = 8'h00; // 0x73e
	13'h73f: qq = 8'h00; // 0x73f
	13'h740: qq = 8'h00; // 0x740
	13'h741: qq = 8'h00; // 0x741
	13'h742: qq = 8'h00; // 0x742
	13'h743: qq = 8'h00; // 0x743
	13'h744: qq = 8'h00; // 0x744
	13'h745: qq = 8'h00; // 0x745
	13'h746: qq = 8'h00; // 0x746
	13'h747: qq = 8'h00; // 0x747
	13'h748: qq = 8'h00; // 0x748
	13'h749: qq = 8'h00; // 0x749
	13'h74a: qq = 8'h00; // 0x74a
	13'h74b: qq = 8'h00; // 0x74b
	13'h74c: qq = 8'h00; // 0x74c
	13'h74d: qq = 8'h00; // 0x74d
	13'h74e: qq = 8'h00; // 0x74e
	13'h74f: qq = 8'h00; // 0x74f
	13'h750: qq = 8'h00; // 0x750
	13'h751: qq = 8'h00; // 0x751
	13'h752: qq = 8'h00; // 0x752
	13'h753: qq = 8'h00; // 0x753
	13'h754: qq = 8'h00; // 0x754
	13'h755: qq = 8'h00; // 0x755
	13'h756: qq = 8'h00; // 0x756
	13'h757: qq = 8'h00; // 0x757
	13'h758: qq = 8'h00; // 0x758
	13'h759: qq = 8'h00; // 0x759
	13'h75a: qq = 8'h00; // 0x75a
	13'h75b: qq = 8'h00; // 0x75b
	13'h75c: qq = 8'h00; // 0x75c
	13'h75d: qq = 8'h00; // 0x75d
	13'h75e: qq = 8'h00; // 0x75e
	13'h75f: qq = 8'h00; // 0x75f
	13'h760: qq = 8'h00; // 0x760
	13'h761: qq = 8'h00; // 0x761
	13'h762: qq = 8'h00; // 0x762
	13'h763: qq = 8'h00; // 0x763
	13'h764: qq = 8'h00; // 0x764
	13'h765: qq = 8'h00; // 0x765
	13'h766: qq = 8'h00; // 0x766
	13'h767: qq = 8'h00; // 0x767
	13'h768: qq = 8'h00; // 0x768
	13'h769: qq = 8'h00; // 0x769
	13'h76a: qq = 8'h00; // 0x76a
	13'h76b: qq = 8'h00; // 0x76b
	13'h76c: qq = 8'h00; // 0x76c
	13'h76d: qq = 8'h00; // 0x76d
	13'h76e: qq = 8'h00; // 0x76e
	13'h76f: qq = 8'h00; // 0x76f
	13'h770: qq = 8'h00; // 0x770
	13'h771: qq = 8'h00; // 0x771
	13'h772: qq = 8'h00; // 0x772
	13'h773: qq = 8'h00; // 0x773
	13'h774: qq = 8'h00; // 0x774
	13'h775: qq = 8'h00; // 0x775
	13'h776: qq = 8'h00; // 0x776
	13'h777: qq = 8'h00; // 0x777
	13'h778: qq = 8'h00; // 0x778
	13'h779: qq = 8'h00; // 0x779
	13'h77a: qq = 8'h00; // 0x77a
	13'h77b: qq = 8'h00; // 0x77b
	13'h77c: qq = 8'h00; // 0x77c
	13'h77d: qq = 8'h00; // 0x77d
	13'h77e: qq = 8'h00; // 0x77e
	13'h77f: qq = 8'h00; // 0x77f
	13'h780: qq = 8'h00; // 0x780
	13'h781: qq = 8'h00; // 0x781
	13'h782: qq = 8'h00; // 0x782
	13'h783: qq = 8'h00; // 0x783
	13'h784: qq = 8'h00; // 0x784
	13'h785: qq = 8'h00; // 0x785
	13'h786: qq = 8'h00; // 0x786
	13'h787: qq = 8'h00; // 0x787
	13'h788: qq = 8'h00; // 0x788
	13'h789: qq = 8'h00; // 0x789
	13'h78a: qq = 8'h00; // 0x78a
	13'h78b: qq = 8'h00; // 0x78b
	13'h78c: qq = 8'h00; // 0x78c
	13'h78d: qq = 8'h00; // 0x78d
	13'h78e: qq = 8'h00; // 0x78e
	13'h78f: qq = 8'h00; // 0x78f
	13'h790: qq = 8'h00; // 0x790
	13'h791: qq = 8'h00; // 0x791
	13'h792: qq = 8'h00; // 0x792
	13'h793: qq = 8'h00; // 0x793
	13'h794: qq = 8'h00; // 0x794
	13'h795: qq = 8'h00; // 0x795
	13'h796: qq = 8'h00; // 0x796
	13'h797: qq = 8'h00; // 0x797
	13'h798: qq = 8'h00; // 0x798
	13'h799: qq = 8'h00; // 0x799
	13'h79a: qq = 8'h00; // 0x79a
	13'h79b: qq = 8'h00; // 0x79b
	13'h79c: qq = 8'h00; // 0x79c
	13'h79d: qq = 8'h00; // 0x79d
	13'h79e: qq = 8'h00; // 0x79e
	13'h79f: qq = 8'h00; // 0x79f
	13'h7a0: qq = 8'h00; // 0x7a0
	13'h7a1: qq = 8'h00; // 0x7a1
	13'h7a2: qq = 8'h00; // 0x7a2
	13'h7a3: qq = 8'h00; // 0x7a3
	13'h7a4: qq = 8'h00; // 0x7a4
	13'h7a5: qq = 8'h00; // 0x7a5
	13'h7a6: qq = 8'h00; // 0x7a6
	13'h7a7: qq = 8'h00; // 0x7a7
	13'h7a8: qq = 8'h00; // 0x7a8
	13'h7a9: qq = 8'h00; // 0x7a9
	13'h7aa: qq = 8'h00; // 0x7aa
	13'h7ab: qq = 8'h00; // 0x7ab
	13'h7ac: qq = 8'h00; // 0x7ac
	13'h7ad: qq = 8'h00; // 0x7ad
	13'h7ae: qq = 8'h00; // 0x7ae
	13'h7af: qq = 8'h00; // 0x7af
	13'h7b0: qq = 8'h00; // 0x7b0
	13'h7b1: qq = 8'h00; // 0x7b1
	13'h7b2: qq = 8'h00; // 0x7b2
	13'h7b3: qq = 8'h00; // 0x7b3
	13'h7b4: qq = 8'h00; // 0x7b4
	13'h7b5: qq = 8'h00; // 0x7b5
	13'h7b6: qq = 8'h00; // 0x7b6
	13'h7b7: qq = 8'h00; // 0x7b7
	13'h7b8: qq = 8'h00; // 0x7b8
	13'h7b9: qq = 8'h00; // 0x7b9
	13'h7ba: qq = 8'h00; // 0x7ba
	13'h7bb: qq = 8'h00; // 0x7bb
	13'h7bc: qq = 8'h00; // 0x7bc
	13'h7bd: qq = 8'h00; // 0x7bd
	13'h7be: qq = 8'h00; // 0x7be
	13'h7bf: qq = 8'h00; // 0x7bf
	13'h7c0: qq = 8'h00; // 0x7c0
	13'h7c1: qq = 8'h00; // 0x7c1
	13'h7c2: qq = 8'h00; // 0x7c2
	13'h7c3: qq = 8'h00; // 0x7c3
	13'h7c4: qq = 8'h00; // 0x7c4
	13'h7c5: qq = 8'h00; // 0x7c5
	13'h7c6: qq = 8'h00; // 0x7c6
	13'h7c7: qq = 8'h00; // 0x7c7
	13'h7c8: qq = 8'h00; // 0x7c8
	13'h7c9: qq = 8'h00; // 0x7c9
	13'h7ca: qq = 8'h00; // 0x7ca
	13'h7cb: qq = 8'h00; // 0x7cb
	13'h7cc: qq = 8'h00; // 0x7cc
	13'h7cd: qq = 8'h00; // 0x7cd
	13'h7ce: qq = 8'h00; // 0x7ce
	13'h7cf: qq = 8'h00; // 0x7cf
	13'h7d0: qq = 8'h00; // 0x7d0
	13'h7d1: qq = 8'h00; // 0x7d1
	13'h7d2: qq = 8'h00; // 0x7d2
	13'h7d3: qq = 8'h00; // 0x7d3
	13'h7d4: qq = 8'h00; // 0x7d4
	13'h7d5: qq = 8'h00; // 0x7d5
	13'h7d6: qq = 8'h00; // 0x7d6
	13'h7d7: qq = 8'h00; // 0x7d7
	13'h7d8: qq = 8'h00; // 0x7d8
	13'h7d9: qq = 8'h00; // 0x7d9
	13'h7da: qq = 8'h00; // 0x7da
	13'h7db: qq = 8'h00; // 0x7db
	13'h7dc: qq = 8'h00; // 0x7dc
	13'h7dd: qq = 8'h00; // 0x7dd
	13'h7de: qq = 8'h00; // 0x7de
	13'h7df: qq = 8'h00; // 0x7df
	13'h7e0: qq = 8'h00; // 0x7e0
	13'h7e1: qq = 8'h00; // 0x7e1
	13'h7e2: qq = 8'h00; // 0x7e2
	13'h7e3: qq = 8'h00; // 0x7e3
	13'h7e4: qq = 8'h00; // 0x7e4
	13'h7e5: qq = 8'h00; // 0x7e5
	13'h7e6: qq = 8'h00; // 0x7e6
	13'h7e7: qq = 8'h00; // 0x7e7
	13'h7e8: qq = 8'h00; // 0x7e8
	13'h7e9: qq = 8'h00; // 0x7e9
	13'h7ea: qq = 8'h00; // 0x7ea
	13'h7eb: qq = 8'h00; // 0x7eb
	13'h7ec: qq = 8'h00; // 0x7ec
	13'h7ed: qq = 8'h00; // 0x7ed
	13'h7ee: qq = 8'h00; // 0x7ee
	13'h7ef: qq = 8'h00; // 0x7ef
	13'h7f0: qq = 8'h00; // 0x7f0
	13'h7f1: qq = 8'h00; // 0x7f1
	13'h7f2: qq = 8'h00; // 0x7f2
	13'h7f3: qq = 8'h00; // 0x7f3
	13'h7f4: qq = 8'h00; // 0x7f4
	13'h7f5: qq = 8'h00; // 0x7f5
	13'h7f6: qq = 8'h00; // 0x7f6
	13'h7f7: qq = 8'h00; // 0x7f7
	13'h7f8: qq = 8'h00; // 0x7f8
	13'h7f9: qq = 8'h00; // 0x7f9
	13'h7fa: qq = 8'h00; // 0x7fa
	13'h7fb: qq = 8'h30; // 0x7fb
	13'h7fc: qq = 8'h3c; // 0x7fc
	13'h7fd: qq = 8'h30; // 0x7fd
	13'h7fe: qq = 8'h3c; // 0x7fe
	13'h7ff: qq = 8'h30; // 0x7ff
		endcase

	assign q = qq;
	endmodule // rom prog_rom4
