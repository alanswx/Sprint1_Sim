library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
ENTITY sync_prom IS
PORT
(
	address         : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	clock           : IN STD_LOGIC  := '1';
	q               : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
);
END sync_prom; 
ARCHITECTURE SYN OF sync_prom IS	
signal qq : STD_LOGIC_VECTOR (3 DOWNTO 0);
begin
q<=qq;
PROCESS (address)
begin
CASE address IS 
	when "00000000" => qq <= "0000"; -- 0x000
	when "00000001" => qq <= "0000"; -- 0x001
	when "00000010" => qq <= "0000"; -- 0x002
	when "00000011" => qq <= "0000"; -- 0x003
	when "00000100" => qq <= "0000"; -- 0x004
	when "00000101" => qq <= "0000"; -- 0x005
	when "00000110" => qq <= "0000"; -- 0x006
	when "00000111" => qq <= "0000"; -- 0x007
	when "00001000" => qq <= "0000"; -- 0x008
	when "00001001" => qq <= "0000"; -- 0x009
	when "00001010" => qq <= "0000"; -- 0x00a
	when "00001011" => qq <= "0000"; -- 0x00b
	when "00001100" => qq <= "0000"; -- 0x00c
	when "00001101" => qq <= "0000"; -- 0x00d
	when "00001110" => qq <= "0000"; -- 0x00e
	when "00001111" => qq <= "0000"; -- 0x00f
	when "00010000" => qq <= "0000"; -- 0x010
	when "00010001" => qq <= "0000"; -- 0x011
	when "00010010" => qq <= "0000"; -- 0x012
	when "00010011" => qq <= "0000"; -- 0x013
	when "00010100" => qq <= "0000"; -- 0x014
	when "00010101" => qq <= "0000"; -- 0x015
	when "00010110" => qq <= "0000"; -- 0x016
	when "00010111" => qq <= "0000"; -- 0x017
	when "00011000" => qq <= "0000"; -- 0x018
	when "00011001" => qq <= "0000"; -- 0x019
	when "00011010" => qq <= "0000"; -- 0x01a
	when "00011011" => qq <= "0000"; -- 0x01b
	when "00011100" => qq <= "0000"; -- 0x01c
	when "00011101" => qq <= "0000"; -- 0x01d
	when "00011110" => qq <= "0000"; -- 0x01e
	when "00011111" => qq <= "0000"; -- 0x01f
	when "00100000" => qq <= "0000"; -- 0x020
	when "00100001" => qq <= "0000"; -- 0x021
	when "00100010" => qq <= "0000"; -- 0x022
	when "00100011" => qq <= "0000"; -- 0x023
	when "00100100" => qq <= "0000"; -- 0x024
	when "00100101" => qq <= "0000"; -- 0x025
	when "00100110" => qq <= "0000"; -- 0x026
	when "00100111" => qq <= "0000"; -- 0x027
	when "00101000" => qq <= "0000"; -- 0x028
	when "00101001" => qq <= "0000"; -- 0x029
	when "00101010" => qq <= "0000"; -- 0x02a
	when "00101011" => qq <= "0000"; -- 0x02b
	when "00101100" => qq <= "0000"; -- 0x02c
	when "00101101" => qq <= "0000"; -- 0x02d
	when "00101110" => qq <= "0000"; -- 0x02e
	when "00101111" => qq <= "0000"; -- 0x02f
	when "00110000" => qq <= "0000"; -- 0x030
	when "00110001" => qq <= "0000"; -- 0x031
	when "00110010" => qq <= "0000"; -- 0x032
	when "00110011" => qq <= "0000"; -- 0x033
	when "00110100" => qq <= "0000"; -- 0x034
	when "00110101" => qq <= "0000"; -- 0x035
	when "00110110" => qq <= "0000"; -- 0x036
	when "00110111" => qq <= "0000"; -- 0x037
	when "00111000" => qq <= "0000"; -- 0x038
	when "00111001" => qq <= "0000"; -- 0x039
	when "00111010" => qq <= "0000"; -- 0x03a
	when "00111011" => qq <= "0000"; -- 0x03b
	when "00111100" => qq <= "0000"; -- 0x03c
	when "00111101" => qq <= "0000"; -- 0x03d
	when "00111110" => qq <= "0000"; -- 0x03e
	when "00111111" => qq <= "0000"; -- 0x03f
	when "01000000" => qq <= "0000"; -- 0x040
	when "01000001" => qq <= "0000"; -- 0x041
	when "01000010" => qq <= "0000"; -- 0x042
	when "01000011" => qq <= "0000"; -- 0x043
	when "01000100" => qq <= "0000"; -- 0x044
	when "01000101" => qq <= "0000"; -- 0x045
	when "01000110" => qq <= "0000"; -- 0x046
	when "01000111" => qq <= "0000"; -- 0x047
	when "01001000" => qq <= "0000"; -- 0x048
	when "01001001" => qq <= "0000"; -- 0x049
	when "01001010" => qq <= "0000"; -- 0x04a
	when "01001011" => qq <= "0000"; -- 0x04b
	when "01001100" => qq <= "0000"; -- 0x04c
	when "01001101" => qq <= "0000"; -- 0x04d
	when "01001110" => qq <= "0000"; -- 0x04e
	when "01001111" => qq <= "0000"; -- 0x04f
	when "01010000" => qq <= "0000"; -- 0x050
	when "01010001" => qq <= "0000"; -- 0x051
	when "01010010" => qq <= "0000"; -- 0x052
	when "01010011" => qq <= "0000"; -- 0x053
	when "01010100" => qq <= "0000"; -- 0x054
	when "01010101" => qq <= "0000"; -- 0x055
	when "01010110" => qq <= "0000"; -- 0x056
	when "01010111" => qq <= "0000"; -- 0x057
	when "01011000" => qq <= "0000"; -- 0x058
	when "01011001" => qq <= "0000"; -- 0x059
	when "01011010" => qq <= "0000"; -- 0x05a
	when "01011011" => qq <= "0000"; -- 0x05b
	when "01011100" => qq <= "0000"; -- 0x05c
	when "01011101" => qq <= "0000"; -- 0x05d
	when "01011110" => qq <= "0000"; -- 0x05e
	when "01011111" => qq <= "0000"; -- 0x05f
	when "01100000" => qq <= "0000"; -- 0x060
	when "01100001" => qq <= "0000"; -- 0x061
	when "01100010" => qq <= "0000"; -- 0x062
	when "01100011" => qq <= "0000"; -- 0x063
	when "01100100" => qq <= "0000"; -- 0x064
	when "01100101" => qq <= "0000"; -- 0x065
	when "01100110" => qq <= "0000"; -- 0x066
	when "01100111" => qq <= "0000"; -- 0x067
	when "01101000" => qq <= "0000"; -- 0x068
	when "01101001" => qq <= "0000"; -- 0x069
	when "01101010" => qq <= "0000"; -- 0x06a
	when "01101011" => qq <= "0000"; -- 0x06b
	when "01101100" => qq <= "0000"; -- 0x06c
	when "01101101" => qq <= "0000"; -- 0x06d
	when "01101110" => qq <= "0000"; -- 0x06e
	when "01101111" => qq <= "0000"; -- 0x06f
	when "01110000" => qq <= "0000"; -- 0x070
	when "01110001" => qq <= "0000"; -- 0x071
	when "01110010" => qq <= "0000"; -- 0x072
	when "01110011" => qq <= "0000"; -- 0x073
	when "01110100" => qq <= "0000"; -- 0x074
	when "01110101" => qq <= "0000"; -- 0x075
	when "01110110" => qq <= "0000"; -- 0x076
	when "01110111" => qq <= "0000"; -- 0x077
	when "01111000" => qq <= "0000"; -- 0x078
	when "01111001" => qq <= "0000"; -- 0x079
	when "01111010" => qq <= "0000"; -- 0x07a
	when "01111011" => qq <= "0000"; -- 0x07b
	when "01111100" => qq <= "0000"; -- 0x07c
	when "01111101" => qq <= "0000"; -- 0x07d
	when "01111110" => qq <= "0000"; -- 0x07e
	when "01111111" => qq <= "1000"; -- 0x07f
	when "10000000" => qq <= "1010"; -- 0x080
	when "10000001" => qq <= "1010"; -- 0x081
	when "10000010" => qq <= "1010"; -- 0x082
	when "10000011" => qq <= "1010"; -- 0x083
	when "10000100" => qq <= "1010"; -- 0x084
	when "10000101" => qq <= "1110"; -- 0x085
	when "10000110" => qq <= "0000"; -- 0x086
	when "10000111" => qq <= "0000"; -- 0x087
	when "10001000" => qq <= "0000"; -- 0x088
	when "10001001" => qq <= "0000"; -- 0x089
	when "10001010" => qq <= "0000"; -- 0x08a
	when "10001011" => qq <= "0000"; -- 0x08b
	when "10001100" => qq <= "0000"; -- 0x08c
	when "10001101" => qq <= "0000"; -- 0x08d
	when "10001110" => qq <= "0000"; -- 0x08e
	when "10001111" => qq <= "0000"; -- 0x08f
	when "10010000" => qq <= "0000"; -- 0x090
	when "10010001" => qq <= "0000"; -- 0x091
	when "10010010" => qq <= "0000"; -- 0x092
	when "10010011" => qq <= "0000"; -- 0x093
	when "10010100" => qq <= "0000"; -- 0x094
	when "10010101" => qq <= "0000"; -- 0x095
	when "10010110" => qq <= "0000"; -- 0x096
	when "10010111" => qq <= "0000"; -- 0x097
	when "10011000" => qq <= "0000"; -- 0x098
	when "10011001" => qq <= "0000"; -- 0x099
	when "10011010" => qq <= "0000"; -- 0x09a
	when "10011011" => qq <= "0000"; -- 0x09b
	when "10011100" => qq <= "0000"; -- 0x09c
	when "10011101" => qq <= "0000"; -- 0x09d
	when "10011110" => qq <= "0000"; -- 0x09e
	when "10011111" => qq <= "0000"; -- 0x09f
	when "10100000" => qq <= "0000"; -- 0x0a0
	when "10100001" => qq <= "0000"; -- 0x0a1
	when "10100010" => qq <= "0000"; -- 0x0a2
	when "10100011" => qq <= "0000"; -- 0x0a3
	when "10100100" => qq <= "0000"; -- 0x0a4
	when "10100101" => qq <= "0000"; -- 0x0a5
	when "10100110" => qq <= "0000"; -- 0x0a6
	when "10100111" => qq <= "0000"; -- 0x0a7
	when "10101000" => qq <= "0000"; -- 0x0a8
	when "10101001" => qq <= "0000"; -- 0x0a9
	when "10101010" => qq <= "0000"; -- 0x0aa
	when "10101011" => qq <= "0000"; -- 0x0ab
	when "10101100" => qq <= "0000"; -- 0x0ac
	when "10101101" => qq <= "0000"; -- 0x0ad
	when "10101110" => qq <= "0000"; -- 0x0ae
	when "10101111" => qq <= "0000"; -- 0x0af
	when "10110000" => qq <= "0000"; -- 0x0b0
	when "10110001" => qq <= "0000"; -- 0x0b1
	when "10110010" => qq <= "0000"; -- 0x0b2
	when "10110011" => qq <= "0000"; -- 0x0b3
	when "10110100" => qq <= "0000"; -- 0x0b4
	when "10110101" => qq <= "0000"; -- 0x0b5
	when "10110110" => qq <= "0000"; -- 0x0b6
	when "10110111" => qq <= "0000"; -- 0x0b7
	when "10111000" => qq <= "0000"; -- 0x0b8
	when "10111001" => qq <= "0000"; -- 0x0b9
	when "10111010" => qq <= "0000"; -- 0x0ba
	when "10111011" => qq <= "0000"; -- 0x0bb
	when "10111100" => qq <= "0000"; -- 0x0bc
	when "10111101" => qq <= "0000"; -- 0x0bd
	when "10111110" => qq <= "0000"; -- 0x0be
	when "10111111" => qq <= "0000"; -- 0x0bf
	when "11000000" => qq <= "0000"; -- 0x0c0
	when "11000001" => qq <= "0000"; -- 0x0c1
	when "11000010" => qq <= "0000"; -- 0x0c2
	when "11000011" => qq <= "0000"; -- 0x0c3
	when "11000100" => qq <= "0000"; -- 0x0c4
	when "11000101" => qq <= "0000"; -- 0x0c5
	when "11000110" => qq <= "0000"; -- 0x0c6
	when "11000111" => qq <= "0000"; -- 0x0c7
	when "11001000" => qq <= "0000"; -- 0x0c8
	when "11001001" => qq <= "0000"; -- 0x0c9
	when "11001010" => qq <= "0000"; -- 0x0ca
	when "11001011" => qq <= "0000"; -- 0x0cb
	when "11001100" => qq <= "0000"; -- 0x0cc
	when "11001101" => qq <= "0000"; -- 0x0cd
	when "11001110" => qq <= "0000"; -- 0x0ce
	when "11001111" => qq <= "0000"; -- 0x0cf
	when "11010000" => qq <= "0000"; -- 0x0d0
	when "11010001" => qq <= "0000"; -- 0x0d1
	when "11010010" => qq <= "0000"; -- 0x0d2
	when "11010011" => qq <= "0000"; -- 0x0d3
	when "11010100" => qq <= "0000"; -- 0x0d4
	when "11010101" => qq <= "0000"; -- 0x0d5
	when "11010110" => qq <= "0000"; -- 0x0d6
	when "11010111" => qq <= "0000"; -- 0x0d7
	when "11011000" => qq <= "0000"; -- 0x0d8
	when "11011001" => qq <= "0000"; -- 0x0d9
	when "11011010" => qq <= "0000"; -- 0x0da
	when "11011011" => qq <= "0000"; -- 0x0db
	when "11011100" => qq <= "0000"; -- 0x0dc
	when "11011101" => qq <= "0000"; -- 0x0dd
	when "11011110" => qq <= "0000"; -- 0x0de
	when "11011111" => qq <= "0000"; -- 0x0df
	when "11100000" => qq <= "1000"; -- 0x0e0
	when "11100001" => qq <= "1000"; -- 0x0e1
	when "11100010" => qq <= "1000"; -- 0x0e2
	when "11100011" => qq <= "1000"; -- 0x0e3
	when "11100100" => qq <= "1000"; -- 0x0e4
	when "11100101" => qq <= "1000"; -- 0x0e5
	when "11100110" => qq <= "1000"; -- 0x0e6
	when "11100111" => qq <= "1000"; -- 0x0e7
	when "11101000" => qq <= "1000"; -- 0x0e8
	when "11101001" => qq <= "1000"; -- 0x0e9
	when "11101010" => qq <= "1000"; -- 0x0ea
	when "11101011" => qq <= "1000"; -- 0x0eb
	when "11101100" => qq <= "1000"; -- 0x0ec
	when "11101101" => qq <= "1000"; -- 0x0ed
	when "11101110" => qq <= "1000"; -- 0x0ee
	when "11101111" => qq <= "1010"; -- 0x0ef
	when "11110000" => qq <= "1010"; -- 0x0f0
	when "11110001" => qq <= "1010"; -- 0x0f1
	when "11110010" => qq <= "1011"; -- 0x0f2
	when "11110011" => qq <= "1011"; -- 0x0f3
	when "11110100" => qq <= "1011"; -- 0x0f4
	when "11110101" => qq <= "1010"; -- 0x0f5
	when "11110110" => qq <= "1010"; -- 0x0f6
	when "11110111" => qq <= "1010"; -- 0x0f7
	when "11111000" => qq <= "1010"; -- 0x0f8
	when "11111001" => qq <= "1010"; -- 0x0f9
	when "11111010" => qq <= "1010"; -- 0x0fa
	when "11111011" => qq <= "1010"; -- 0x0fb
	when "11111100" => qq <= "1010"; -- 0x0fc
	when "11111101" => qq <= "1010"; -- 0x0fd
	when "11111110" => qq <= "1010"; -- 0x0fe
	when "11111111" => qq <= "1010"; -- 0x0ff
	when others => qq <= "0000";
END CASE; 
END PROCESS; 
END SYN; 
