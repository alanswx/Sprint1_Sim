module sync_prom(input clock,
	input [7:0] address,
	output [3:0] q
	);

	reg [3:0] qq;
always @(posedge clk )
		case (address)
	13'h000: qq = 8'h00; // 0x000
	13'h001: qq = 8'h00; // 0x001
	13'h002: qq = 8'h00; // 0x002
	13'h003: qq = 8'h00; // 0x003
	13'h004: qq = 8'h00; // 0x004
	13'h005: qq = 8'h00; // 0x005
	13'h006: qq = 8'h00; // 0x006
	13'h007: qq = 8'h00; // 0x007
	13'h008: qq = 8'h00; // 0x008
	13'h009: qq = 8'h00; // 0x009
	13'h00a: qq = 8'h00; // 0x00a
	13'h00b: qq = 8'h00; // 0x00b
	13'h00c: qq = 8'h00; // 0x00c
	13'h00d: qq = 8'h00; // 0x00d
	13'h00e: qq = 8'h00; // 0x00e
	13'h00f: qq = 8'h00; // 0x00f
	13'h010: qq = 8'h00; // 0x010
	13'h011: qq = 8'h00; // 0x011
	13'h012: qq = 8'h00; // 0x012
	13'h013: qq = 8'h00; // 0x013
	13'h014: qq = 8'h00; // 0x014
	13'h015: qq = 8'h00; // 0x015
	13'h016: qq = 8'h00; // 0x016
	13'h017: qq = 8'h00; // 0x017
	13'h018: qq = 8'h00; // 0x018
	13'h019: qq = 8'h00; // 0x019
	13'h01a: qq = 8'h00; // 0x01a
	13'h01b: qq = 8'h00; // 0x01b
	13'h01c: qq = 8'h00; // 0x01c
	13'h01d: qq = 8'h00; // 0x01d
	13'h01e: qq = 8'h00; // 0x01e
	13'h01f: qq = 8'h00; // 0x01f
	13'h020: qq = 8'h00; // 0x020
	13'h021: qq = 8'h00; // 0x021
	13'h022: qq = 8'h00; // 0x022
	13'h023: qq = 8'h00; // 0x023
	13'h024: qq = 8'h00; // 0x024
	13'h025: qq = 8'h00; // 0x025
	13'h026: qq = 8'h00; // 0x026
	13'h027: qq = 8'h00; // 0x027
	13'h028: qq = 8'h00; // 0x028
	13'h029: qq = 8'h00; // 0x029
	13'h02a: qq = 8'h00; // 0x02a
	13'h02b: qq = 8'h00; // 0x02b
	13'h02c: qq = 8'h00; // 0x02c
	13'h02d: qq = 8'h00; // 0x02d
	13'h02e: qq = 8'h00; // 0x02e
	13'h02f: qq = 8'h00; // 0x02f
	13'h030: qq = 8'h00; // 0x030
	13'h031: qq = 8'h00; // 0x031
	13'h032: qq = 8'h00; // 0x032
	13'h033: qq = 8'h00; // 0x033
	13'h034: qq = 8'h00; // 0x034
	13'h035: qq = 8'h00; // 0x035
	13'h036: qq = 8'h00; // 0x036
	13'h037: qq = 8'h00; // 0x037
	13'h038: qq = 8'h00; // 0x038
	13'h039: qq = 8'h00; // 0x039
	13'h03a: qq = 8'h00; // 0x03a
	13'h03b: qq = 8'h00; // 0x03b
	13'h03c: qq = 8'h00; // 0x03c
	13'h03d: qq = 8'h00; // 0x03d
	13'h03e: qq = 8'h00; // 0x03e
	13'h03f: qq = 8'h00; // 0x03f
	13'h040: qq = 8'h00; // 0x040
	13'h041: qq = 8'h00; // 0x041
	13'h042: qq = 8'h00; // 0x042
	13'h043: qq = 8'h00; // 0x043
	13'h044: qq = 8'h00; // 0x044
	13'h045: qq = 8'h00; // 0x045
	13'h046: qq = 8'h00; // 0x046
	13'h047: qq = 8'h00; // 0x047
	13'h048: qq = 8'h00; // 0x048
	13'h049: qq = 8'h00; // 0x049
	13'h04a: qq = 8'h00; // 0x04a
	13'h04b: qq = 8'h00; // 0x04b
	13'h04c: qq = 8'h00; // 0x04c
	13'h04d: qq = 8'h00; // 0x04d
	13'h04e: qq = 8'h00; // 0x04e
	13'h04f: qq = 8'h00; // 0x04f
	13'h050: qq = 8'h00; // 0x050
	13'h051: qq = 8'h00; // 0x051
	13'h052: qq = 8'h00; // 0x052
	13'h053: qq = 8'h00; // 0x053
	13'h054: qq = 8'h00; // 0x054
	13'h055: qq = 8'h00; // 0x055
	13'h056: qq = 8'h00; // 0x056
	13'h057: qq = 8'h00; // 0x057
	13'h058: qq = 8'h00; // 0x058
	13'h059: qq = 8'h00; // 0x059
	13'h05a: qq = 8'h00; // 0x05a
	13'h05b: qq = 8'h00; // 0x05b
	13'h05c: qq = 8'h00; // 0x05c
	13'h05d: qq = 8'h00; // 0x05d
	13'h05e: qq = 8'h00; // 0x05e
	13'h05f: qq = 8'h00; // 0x05f
	13'h060: qq = 8'h00; // 0x060
	13'h061: qq = 8'h00; // 0x061
	13'h062: qq = 8'h00; // 0x062
	13'h063: qq = 8'h00; // 0x063
	13'h064: qq = 8'h00; // 0x064
	13'h065: qq = 8'h00; // 0x065
	13'h066: qq = 8'h00; // 0x066
	13'h067: qq = 8'h00; // 0x067
	13'h068: qq = 8'h00; // 0x068
	13'h069: qq = 8'h00; // 0x069
	13'h06a: qq = 8'h00; // 0x06a
	13'h06b: qq = 8'h00; // 0x06b
	13'h06c: qq = 8'h00; // 0x06c
	13'h06d: qq = 8'h00; // 0x06d
	13'h06e: qq = 8'h00; // 0x06e
	13'h06f: qq = 8'h00; // 0x06f
	13'h070: qq = 8'h00; // 0x070
	13'h071: qq = 8'h00; // 0x071
	13'h072: qq = 8'h00; // 0x072
	13'h073: qq = 8'h00; // 0x073
	13'h074: qq = 8'h00; // 0x074
	13'h075: qq = 8'h00; // 0x075
	13'h076: qq = 8'h00; // 0x076
	13'h077: qq = 8'h00; // 0x077
	13'h078: qq = 8'h00; // 0x078
	13'h079: qq = 8'h00; // 0x079
	13'h07a: qq = 8'h00; // 0x07a
	13'h07b: qq = 8'h00; // 0x07b
	13'h07c: qq = 8'h00; // 0x07c
	13'h07d: qq = 8'h00; // 0x07d
	13'h07e: qq = 8'h00; // 0x07e
	13'h07f: qq = 8'h08; // 0x07f
	13'h080: qq = 8'h0a; // 0x080
	13'h081: qq = 8'h0a; // 0x081
	13'h082: qq = 8'h0a; // 0x082
	13'h083: qq = 8'h0a; // 0x083
	13'h084: qq = 8'h0a; // 0x084
	13'h085: qq = 8'h0e; // 0x085
	13'h086: qq = 8'h00; // 0x086
	13'h087: qq = 8'h00; // 0x087
	13'h088: qq = 8'h00; // 0x088
	13'h089: qq = 8'h00; // 0x089
	13'h08a: qq = 8'h00; // 0x08a
	13'h08b: qq = 8'h00; // 0x08b
	13'h08c: qq = 8'h00; // 0x08c
	13'h08d: qq = 8'h00; // 0x08d
	13'h08e: qq = 8'h00; // 0x08e
	13'h08f: qq = 8'h00; // 0x08f
	13'h090: qq = 8'h00; // 0x090
	13'h091: qq = 8'h00; // 0x091
	13'h092: qq = 8'h00; // 0x092
	13'h093: qq = 8'h00; // 0x093
	13'h094: qq = 8'h00; // 0x094
	13'h095: qq = 8'h00; // 0x095
	13'h096: qq = 8'h00; // 0x096
	13'h097: qq = 8'h00; // 0x097
	13'h098: qq = 8'h00; // 0x098
	13'h099: qq = 8'h00; // 0x099
	13'h09a: qq = 8'h00; // 0x09a
	13'h09b: qq = 8'h00; // 0x09b
	13'h09c: qq = 8'h00; // 0x09c
	13'h09d: qq = 8'h00; // 0x09d
	13'h09e: qq = 8'h00; // 0x09e
	13'h09f: qq = 8'h00; // 0x09f
	13'h0a0: qq = 8'h00; // 0x0a0
	13'h0a1: qq = 8'h00; // 0x0a1
	13'h0a2: qq = 8'h00; // 0x0a2
	13'h0a3: qq = 8'h00; // 0x0a3
	13'h0a4: qq = 8'h00; // 0x0a4
	13'h0a5: qq = 8'h00; // 0x0a5
	13'h0a6: qq = 8'h00; // 0x0a6
	13'h0a7: qq = 8'h00; // 0x0a7
	13'h0a8: qq = 8'h00; // 0x0a8
	13'h0a9: qq = 8'h00; // 0x0a9
	13'h0aa: qq = 8'h00; // 0x0aa
	13'h0ab: qq = 8'h00; // 0x0ab
	13'h0ac: qq = 8'h00; // 0x0ac
	13'h0ad: qq = 8'h00; // 0x0ad
	13'h0ae: qq = 8'h00; // 0x0ae
	13'h0af: qq = 8'h00; // 0x0af
	13'h0b0: qq = 8'h00; // 0x0b0
	13'h0b1: qq = 8'h00; // 0x0b1
	13'h0b2: qq = 8'h00; // 0x0b2
	13'h0b3: qq = 8'h00; // 0x0b3
	13'h0b4: qq = 8'h00; // 0x0b4
	13'h0b5: qq = 8'h00; // 0x0b5
	13'h0b6: qq = 8'h00; // 0x0b6
	13'h0b7: qq = 8'h00; // 0x0b7
	13'h0b8: qq = 8'h00; // 0x0b8
	13'h0b9: qq = 8'h00; // 0x0b9
	13'h0ba: qq = 8'h00; // 0x0ba
	13'h0bb: qq = 8'h00; // 0x0bb
	13'h0bc: qq = 8'h00; // 0x0bc
	13'h0bd: qq = 8'h00; // 0x0bd
	13'h0be: qq = 8'h00; // 0x0be
	13'h0bf: qq = 8'h00; // 0x0bf
	13'h0c0: qq = 8'h00; // 0x0c0
	13'h0c1: qq = 8'h00; // 0x0c1
	13'h0c2: qq = 8'h00; // 0x0c2
	13'h0c3: qq = 8'h00; // 0x0c3
	13'h0c4: qq = 8'h00; // 0x0c4
	13'h0c5: qq = 8'h00; // 0x0c5
	13'h0c6: qq = 8'h00; // 0x0c6
	13'h0c7: qq = 8'h00; // 0x0c7
	13'h0c8: qq = 8'h00; // 0x0c8
	13'h0c9: qq = 8'h00; // 0x0c9
	13'h0ca: qq = 8'h00; // 0x0ca
	13'h0cb: qq = 8'h00; // 0x0cb
	13'h0cc: qq = 8'h00; // 0x0cc
	13'h0cd: qq = 8'h00; // 0x0cd
	13'h0ce: qq = 8'h00; // 0x0ce
	13'h0cf: qq = 8'h00; // 0x0cf
	13'h0d0: qq = 8'h00; // 0x0d0
	13'h0d1: qq = 8'h00; // 0x0d1
	13'h0d2: qq = 8'h00; // 0x0d2
	13'h0d3: qq = 8'h00; // 0x0d3
	13'h0d4: qq = 8'h00; // 0x0d4
	13'h0d5: qq = 8'h00; // 0x0d5
	13'h0d6: qq = 8'h00; // 0x0d6
	13'h0d7: qq = 8'h00; // 0x0d7
	13'h0d8: qq = 8'h00; // 0x0d8
	13'h0d9: qq = 8'h00; // 0x0d9
	13'h0da: qq = 8'h00; // 0x0da
	13'h0db: qq = 8'h00; // 0x0db
	13'h0dc: qq = 8'h00; // 0x0dc
	13'h0dd: qq = 8'h00; // 0x0dd
	13'h0de: qq = 8'h00; // 0x0de
	13'h0df: qq = 8'h00; // 0x0df
	13'h0e0: qq = 8'h08; // 0x0e0
	13'h0e1: qq = 8'h08; // 0x0e1
	13'h0e2: qq = 8'h08; // 0x0e2
	13'h0e3: qq = 8'h08; // 0x0e3
	13'h0e4: qq = 8'h08; // 0x0e4
	13'h0e5: qq = 8'h08; // 0x0e5
	13'h0e6: qq = 8'h08; // 0x0e6
	13'h0e7: qq = 8'h08; // 0x0e7
	13'h0e8: qq = 8'h08; // 0x0e8
	13'h0e9: qq = 8'h08; // 0x0e9
	13'h0ea: qq = 8'h08; // 0x0ea
	13'h0eb: qq = 8'h08; // 0x0eb
	13'h0ec: qq = 8'h08; // 0x0ec
	13'h0ed: qq = 8'h08; // 0x0ed
	13'h0ee: qq = 8'h08; // 0x0ee
	13'h0ef: qq = 8'h0a; // 0x0ef
	13'h0f0: qq = 8'h0a; // 0x0f0
	13'h0f1: qq = 8'h0a; // 0x0f1
	13'h0f2: qq = 8'h0b; // 0x0f2
	13'h0f3: qq = 8'h0b; // 0x0f3
	13'h0f4: qq = 8'h0b; // 0x0f4
	13'h0f5: qq = 8'h0a; // 0x0f5
	13'h0f6: qq = 8'h0a; // 0x0f6
	13'h0f7: qq = 8'h0a; // 0x0f7
	13'h0f8: qq = 8'h0a; // 0x0f8
	13'h0f9: qq = 8'h0a; // 0x0f9
	13'h0fa: qq = 8'h0a; // 0x0fa
	13'h0fb: qq = 8'h0a; // 0x0fb
	13'h0fc: qq = 8'h0a; // 0x0fc
	13'h0fd: qq = 8'h0a; // 0x0fd
	13'h0fe: qq = 8'h0a; // 0x0fe
	13'h0ff: qq = 8'h0a; // 0x0ff
		endcase

	assign q = qq;
	endmodule // rom sync_prom
