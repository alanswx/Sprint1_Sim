module Char_MSB(input clock,
	input [8:0] address,
	output [3:0] q
	);

	reg [3:0] qq;
always @(posedge clk )
		case (address)
	13'h000: qq = 8'h00; // 0x000
	13'h001: qq = 8'h00; // 0x001
	13'h002: qq = 8'h00; // 0x002
	13'h003: qq = 8'h00; // 0x003
	13'h004: qq = 8'h00; // 0x004
	13'h005: qq = 8'h00; // 0x005
	13'h006: qq = 8'h00; // 0x006
	13'h007: qq = 8'h00; // 0x007
	13'h008: qq = 8'h00; // 0x008
	13'h009: qq = 8'h08; // 0x009
	13'h00a: qq = 8'h0c; // 0x00a
	13'h00b: qq = 8'h06; // 0x00b
	13'h00c: qq = 8'h06; // 0x00c
	13'h00d: qq = 8'h0e; // 0x00d
	13'h00e: qq = 8'h06; // 0x00e
	13'h00f: qq = 8'h06; // 0x00f
	13'h010: qq = 8'h00; // 0x010
	13'h011: qq = 8'h0c; // 0x011
	13'h012: qq = 8'h06; // 0x012
	13'h013: qq = 8'h06; // 0x013
	13'h014: qq = 8'h0c; // 0x014
	13'h015: qq = 8'h06; // 0x015
	13'h016: qq = 8'h06; // 0x016
	13'h017: qq = 8'h0c; // 0x017
	13'h018: qq = 8'h00; // 0x018
	13'h019: qq = 8'h0c; // 0x019
	13'h01a: qq = 8'h06; // 0x01a
	13'h01b: qq = 8'h00; // 0x01b
	13'h01c: qq = 8'h00; // 0x01c
	13'h01d: qq = 8'h00; // 0x01d
	13'h01e: qq = 8'h06; // 0x01e
	13'h01f: qq = 8'h0c; // 0x01f
	13'h020: qq = 8'h00; // 0x020
	13'h021: qq = 8'h08; // 0x021
	13'h022: qq = 8'h0c; // 0x022
	13'h023: qq = 8'h06; // 0x023
	13'h024: qq = 8'h06; // 0x024
	13'h025: qq = 8'h06; // 0x025
	13'h026: qq = 8'h0c; // 0x026
	13'h027: qq = 8'h08; // 0x027
	13'h028: qq = 8'h00; // 0x028
	13'h029: qq = 8'h0c; // 0x029
	13'h02a: qq = 8'h00; // 0x02a
	13'h02b: qq = 8'h00; // 0x02b
	13'h02c: qq = 8'h08; // 0x02c
	13'h02d: qq = 8'h00; // 0x02d
	13'h02e: qq = 8'h00; // 0x02e
	13'h02f: qq = 8'h0e; // 0x02f
	13'h030: qq = 8'h00; // 0x030
	13'h031: qq = 8'h0e; // 0x031
	13'h032: qq = 8'h00; // 0x032
	13'h033: qq = 8'h00; // 0x033
	13'h034: qq = 8'h0c; // 0x034
	13'h035: qq = 8'h00; // 0x035
	13'h036: qq = 8'h00; // 0x036
	13'h037: qq = 8'h00; // 0x037
	13'h038: qq = 8'h00; // 0x038
	13'h039: qq = 8'h0e; // 0x039
	13'h03a: qq = 8'h00; // 0x03a
	13'h03b: qq = 8'h00; // 0x03b
	13'h03c: qq = 8'h0e; // 0x03c
	13'h03d: qq = 8'h06; // 0x03d
	13'h03e: qq = 8'h06; // 0x03e
	13'h03f: qq = 8'h0e; // 0x03f
	13'h040: qq = 8'h00; // 0x040
	13'h041: qq = 8'h06; // 0x041
	13'h042: qq = 8'h06; // 0x042
	13'h043: qq = 8'h06; // 0x043
	13'h044: qq = 8'h0e; // 0x044
	13'h045: qq = 8'h06; // 0x045
	13'h046: qq = 8'h06; // 0x046
	13'h047: qq = 8'h06; // 0x047
	13'h048: qq = 8'h00; // 0x048
	13'h049: qq = 8'h0c; // 0x049
	13'h04a: qq = 8'h00; // 0x04a
	13'h04b: qq = 8'h00; // 0x04b
	13'h04c: qq = 8'h00; // 0x04c
	13'h04d: qq = 8'h00; // 0x04d
	13'h04e: qq = 8'h00; // 0x04e
	13'h04f: qq = 8'h0c; // 0x04f
	13'h050: qq = 8'h00; // 0x050
	13'h051: qq = 8'h06; // 0x051
	13'h052: qq = 8'h06; // 0x052
	13'h053: qq = 8'h06; // 0x053
	13'h054: qq = 8'h06; // 0x054
	13'h055: qq = 8'h06; // 0x055
	13'h056: qq = 8'h06; // 0x056
	13'h057: qq = 8'h0c; // 0x057
	13'h058: qq = 8'h00; // 0x058
	13'h059: qq = 8'h06; // 0x059
	13'h05a: qq = 8'h0c; // 0x05a
	13'h05b: qq = 8'h08; // 0x05b
	13'h05c: qq = 8'h00; // 0x05c
	13'h05d: qq = 8'h08; // 0x05d
	13'h05e: qq = 8'h0c; // 0x05e
	13'h05f: qq = 8'h0e; // 0x05f
	13'h060: qq = 8'h00; // 0x060
	13'h061: qq = 8'h00; // 0x061
	13'h062: qq = 8'h00; // 0x062
	13'h063: qq = 8'h00; // 0x063
	13'h064: qq = 8'h00; // 0x064
	13'h065: qq = 8'h00; // 0x065
	13'h066: qq = 8'h00; // 0x066
	13'h067: qq = 8'h0c; // 0x067
	13'h068: qq = 8'h00; // 0x068
	13'h069: qq = 8'h06; // 0x069
	13'h06a: qq = 8'h0e; // 0x06a
	13'h06b: qq = 8'h0e; // 0x06b
	13'h06c: qq = 8'h0e; // 0x06c
	13'h06d: qq = 8'h06; // 0x06d
	13'h06e: qq = 8'h06; // 0x06e
	13'h06f: qq = 8'h06; // 0x06f
	13'h070: qq = 8'h00; // 0x070
	13'h071: qq = 8'h06; // 0x071
	13'h072: qq = 8'h06; // 0x072
	13'h073: qq = 8'h06; // 0x073
	13'h074: qq = 8'h0e; // 0x074
	13'h075: qq = 8'h0e; // 0x075
	13'h076: qq = 8'h0e; // 0x076
	13'h077: qq = 8'h06; // 0x077
	13'h078: qq = 8'h00; // 0x078
	13'h079: qq = 8'h0c; // 0x079
	13'h07a: qq = 8'h06; // 0x07a
	13'h07b: qq = 8'h06; // 0x07b
	13'h07c: qq = 8'h06; // 0x07c
	13'h07d: qq = 8'h06; // 0x07d
	13'h07e: qq = 8'h06; // 0x07e
	13'h07f: qq = 8'h0c; // 0x07f
	13'h080: qq = 8'h00; // 0x080
	13'h081: qq = 8'h0c; // 0x081
	13'h082: qq = 8'h06; // 0x082
	13'h083: qq = 8'h06; // 0x083
	13'h084: qq = 8'h06; // 0x084
	13'h085: qq = 8'h0c; // 0x085
	13'h086: qq = 8'h00; // 0x086
	13'h087: qq = 8'h00; // 0x087
	13'h088: qq = 8'h00; // 0x088
	13'h089: qq = 8'h0c; // 0x089
	13'h08a: qq = 8'h06; // 0x08a
	13'h08b: qq = 8'h06; // 0x08b
	13'h08c: qq = 8'h06; // 0x08c
	13'h08d: qq = 8'h0e; // 0x08d
	13'h08e: qq = 8'h0c; // 0x08e
	13'h08f: qq = 8'h0a; // 0x08f
	13'h090: qq = 8'h00; // 0x090
	13'h091: qq = 8'h0c; // 0x091
	13'h092: qq = 8'h06; // 0x092
	13'h093: qq = 8'h06; // 0x093
	13'h094: qq = 8'h0e; // 0x094
	13'h095: qq = 8'h08; // 0x095
	13'h096: qq = 8'h0c; // 0x096
	13'h097: qq = 8'h0e; // 0x097
	13'h098: qq = 8'h00; // 0x098
	13'h099: qq = 8'h08; // 0x099
	13'h09a: qq = 8'h0c; // 0x09a
	13'h09b: qq = 8'h00; // 0x09b
	13'h09c: qq = 8'h0c; // 0x09c
	13'h09d: qq = 8'h06; // 0x09d
	13'h09e: qq = 8'h06; // 0x09e
	13'h09f: qq = 8'h0c; // 0x09f
	13'h0a0: qq = 8'h00; // 0x0a0
	13'h0a1: qq = 8'h0c; // 0x0a1
	13'h0a2: qq = 8'h00; // 0x0a2
	13'h0a3: qq = 8'h00; // 0x0a3
	13'h0a4: qq = 8'h00; // 0x0a4
	13'h0a5: qq = 8'h00; // 0x0a5
	13'h0a6: qq = 8'h00; // 0x0a6
	13'h0a7: qq = 8'h00; // 0x0a7
	13'h0a8: qq = 8'h00; // 0x0a8
	13'h0a9: qq = 8'h06; // 0x0a9
	13'h0aa: qq = 8'h06; // 0x0aa
	13'h0ab: qq = 8'h06; // 0x0ab
	13'h0ac: qq = 8'h06; // 0x0ac
	13'h0ad: qq = 8'h06; // 0x0ad
	13'h0ae: qq = 8'h06; // 0x0ae
	13'h0af: qq = 8'h0c; // 0x0af
	13'h0b0: qq = 8'h00; // 0x0b0
	13'h0b1: qq = 8'h06; // 0x0b1
	13'h0b2: qq = 8'h06; // 0x0b2
	13'h0b3: qq = 8'h06; // 0x0b3
	13'h0b4: qq = 8'h0e; // 0x0b4
	13'h0b5: qq = 8'h0c; // 0x0b5
	13'h0b6: qq = 8'h08; // 0x0b6
	13'h0b7: qq = 8'h00; // 0x0b7
	13'h0b8: qq = 8'h00; // 0x0b8
	13'h0b9: qq = 8'h06; // 0x0b9
	13'h0ba: qq = 8'h06; // 0x0ba
	13'h0bb: qq = 8'h06; // 0x0bb
	13'h0bc: qq = 8'h0e; // 0x0bc
	13'h0bd: qq = 8'h0e; // 0x0bd
	13'h0be: qq = 8'h0e; // 0x0be
	13'h0bf: qq = 8'h06; // 0x0bf
	13'h0c0: qq = 8'h00; // 0x0c0
	13'h0c1: qq = 8'h06; // 0x0c1
	13'h0c2: qq = 8'h0e; // 0x0c2
	13'h0c3: qq = 8'h0c; // 0x0c3
	13'h0c4: qq = 8'h08; // 0x0c4
	13'h0c5: qq = 8'h0c; // 0x0c5
	13'h0c6: qq = 8'h0e; // 0x0c6
	13'h0c7: qq = 8'h06; // 0x0c7
	13'h0c8: qq = 8'h00; // 0x0c8
	13'h0c9: qq = 8'h0c; // 0x0c9
	13'h0ca: qq = 8'h0c; // 0x0ca
	13'h0cb: qq = 8'h0c; // 0x0cb
	13'h0cc: qq = 8'h08; // 0x0cc
	13'h0cd: qq = 8'h00; // 0x0cd
	13'h0ce: qq = 8'h00; // 0x0ce
	13'h0cf: qq = 8'h00; // 0x0cf
	13'h0d0: qq = 8'h00; // 0x0d0
	13'h0d1: qq = 8'h0e; // 0x0d1
	13'h0d2: qq = 8'h0e; // 0x0d2
	13'h0d3: qq = 8'h0c; // 0x0d3
	13'h0d4: qq = 8'h08; // 0x0d4
	13'h0d5: qq = 8'h00; // 0x0d5
	13'h0d6: qq = 8'h00; // 0x0d6
	13'h0d7: qq = 8'h0e; // 0x0d7
	13'h0d8: qq = 8'h00; // 0x0d8
	13'h0d9: qq = 8'h00; // 0x0d9
	13'h0da: qq = 8'h00; // 0x0da
	13'h0db: qq = 8'h00; // 0x0db
	13'h0dc: qq = 8'h00; // 0x0dc
	13'h0dd: qq = 8'h00; // 0x0dd
	13'h0de: qq = 8'h00; // 0x0de
	13'h0df: qq = 8'h00; // 0x0df
	13'h0e0: qq = 8'h00; // 0x0e0
	13'h0e1: qq = 8'h00; // 0x0e1
	13'h0e2: qq = 8'h00; // 0x0e2
	13'h0e3: qq = 8'h00; // 0x0e3
	13'h0e4: qq = 8'h00; // 0x0e4
	13'h0e5: qq = 8'h00; // 0x0e5
	13'h0e6: qq = 8'h00; // 0x0e6
	13'h0e7: qq = 8'h00; // 0x0e7
	13'h0e8: qq = 8'h00; // 0x0e8
	13'h0e9: qq = 8'h00; // 0x0e9
	13'h0ea: qq = 8'h00; // 0x0ea
	13'h0eb: qq = 8'h00; // 0x0eb
	13'h0ec: qq = 8'h00; // 0x0ec
	13'h0ed: qq = 8'h00; // 0x0ed
	13'h0ee: qq = 8'h00; // 0x0ee
	13'h0ef: qq = 8'h00; // 0x0ef
	13'h0f0: qq = 8'h00; // 0x0f0
	13'h0f1: qq = 8'h00; // 0x0f1
	13'h0f2: qq = 8'h00; // 0x0f2
	13'h0f3: qq = 8'h00; // 0x0f3
	13'h0f4: qq = 8'h00; // 0x0f4
	13'h0f5: qq = 8'h00; // 0x0f5
	13'h0f6: qq = 8'h00; // 0x0f6
	13'h0f7: qq = 8'h00; // 0x0f7
	13'h0f8: qq = 8'h00; // 0x0f8
	13'h0f9: qq = 8'h00; // 0x0f9
	13'h0fa: qq = 8'h00; // 0x0fa
	13'h0fb: qq = 8'h00; // 0x0fb
	13'h0fc: qq = 8'h00; // 0x0fc
	13'h0fd: qq = 8'h00; // 0x0fd
	13'h0fe: qq = 8'h00; // 0x0fe
	13'h0ff: qq = 8'h00; // 0x0ff
	13'h100: qq = 8'h00; // 0x100
	13'h101: qq = 8'h00; // 0x101
	13'h102: qq = 8'h00; // 0x102
	13'h103: qq = 8'h00; // 0x103
	13'h104: qq = 8'h00; // 0x104
	13'h105: qq = 8'h00; // 0x105
	13'h106: qq = 8'h00; // 0x106
	13'h107: qq = 8'h00; // 0x107
	13'h108: qq = 8'h00; // 0x108
	13'h109: qq = 8'h00; // 0x109
	13'h10a: qq = 8'h00; // 0x10a
	13'h10b: qq = 8'h00; // 0x10b
	13'h10c: qq = 8'h00; // 0x10c
	13'h10d: qq = 8'h00; // 0x10d
	13'h10e: qq = 8'h00; // 0x10e
	13'h10f: qq = 8'h00; // 0x10f
	13'h110: qq = 8'h00; // 0x110
	13'h111: qq = 8'h00; // 0x111
	13'h112: qq = 8'h00; // 0x112
	13'h113: qq = 8'h00; // 0x113
	13'h114: qq = 8'h00; // 0x114
	13'h115: qq = 8'h00; // 0x115
	13'h116: qq = 8'h00; // 0x116
	13'h117: qq = 8'h00; // 0x117
	13'h118: qq = 8'h00; // 0x118
	13'h119: qq = 8'h00; // 0x119
	13'h11a: qq = 8'h00; // 0x11a
	13'h11b: qq = 8'h00; // 0x11b
	13'h11c: qq = 8'h00; // 0x11c
	13'h11d: qq = 8'h00; // 0x11d
	13'h11e: qq = 8'h00; // 0x11e
	13'h11f: qq = 8'h00; // 0x11f
	13'h120: qq = 8'h00; // 0x120
	13'h121: qq = 8'h00; // 0x121
	13'h122: qq = 8'h00; // 0x122
	13'h123: qq = 8'h00; // 0x123
	13'h124: qq = 8'h00; // 0x124
	13'h125: qq = 8'h00; // 0x125
	13'h126: qq = 8'h00; // 0x126
	13'h127: qq = 8'h00; // 0x127
	13'h128: qq = 8'h00; // 0x128
	13'h129: qq = 8'h00; // 0x129
	13'h12a: qq = 8'h00; // 0x12a
	13'h12b: qq = 8'h00; // 0x12b
	13'h12c: qq = 8'h00; // 0x12c
	13'h12d: qq = 8'h00; // 0x12d
	13'h12e: qq = 8'h00; // 0x12e
	13'h12f: qq = 8'h00; // 0x12f
	13'h130: qq = 8'h00; // 0x130
	13'h131: qq = 8'h00; // 0x131
	13'h132: qq = 8'h00; // 0x132
	13'h133: qq = 8'h00; // 0x133
	13'h134: qq = 8'h00; // 0x134
	13'h135: qq = 8'h00; // 0x135
	13'h136: qq = 8'h00; // 0x136
	13'h137: qq = 8'h00; // 0x137
	13'h138: qq = 8'h00; // 0x138
	13'h139: qq = 8'h00; // 0x139
	13'h13a: qq = 8'h00; // 0x13a
	13'h13b: qq = 8'h00; // 0x13b
	13'h13c: qq = 8'h00; // 0x13c
	13'h13d: qq = 8'h00; // 0x13d
	13'h13e: qq = 8'h00; // 0x13e
	13'h13f: qq = 8'h00; // 0x13f
	13'h140: qq = 8'h00; // 0x140
	13'h141: qq = 8'h00; // 0x141
	13'h142: qq = 8'h00; // 0x142
	13'h143: qq = 8'h00; // 0x143
	13'h144: qq = 8'h00; // 0x144
	13'h145: qq = 8'h06; // 0x145
	13'h146: qq = 8'h06; // 0x146
	13'h147: qq = 8'h00; // 0x147
	13'h148: qq = 8'h00; // 0x148
	13'h149: qq = 8'h00; // 0x149
	13'h14a: qq = 8'h00; // 0x14a
	13'h14b: qq = 8'h00; // 0x14b
	13'h14c: qq = 8'h00; // 0x14c
	13'h14d: qq = 8'h00; // 0x14d
	13'h14e: qq = 8'h00; // 0x14e
	13'h14f: qq = 8'h00; // 0x14f
	13'h150: qq = 8'h00; // 0x150
	13'h151: qq = 8'h00; // 0x151
	13'h152: qq = 8'h00; // 0x152
	13'h153: qq = 8'h00; // 0x153
	13'h154: qq = 8'h00; // 0x154
	13'h155: qq = 8'h00; // 0x155
	13'h156: qq = 8'h00; // 0x156
	13'h157: qq = 8'h00; // 0x157
	13'h158: qq = 8'h00; // 0x158
	13'h159: qq = 8'h00; // 0x159
	13'h15a: qq = 8'h00; // 0x15a
	13'h15b: qq = 8'h00; // 0x15b
	13'h15c: qq = 8'h00; // 0x15c
	13'h15d: qq = 8'h00; // 0x15d
	13'h15e: qq = 8'h00; // 0x15e
	13'h15f: qq = 8'h00; // 0x15f
	13'h160: qq = 8'h00; // 0x160
	13'h161: qq = 8'h06; // 0x161
	13'h162: qq = 8'h06; // 0x162
	13'h163: qq = 8'h00; // 0x163
	13'h164: qq = 8'h00; // 0x164
	13'h165: qq = 8'h00; // 0x165
	13'h166: qq = 8'h00; // 0x166
	13'h167: qq = 8'h00; // 0x167
	13'h168: qq = 8'h00; // 0x168
	13'h169: qq = 8'h06; // 0x169
	13'h16a: qq = 8'h06; // 0x16a
	13'h16b: qq = 8'h00; // 0x16b
	13'h16c: qq = 8'h00; // 0x16c
	13'h16d: qq = 8'h00; // 0x16d
	13'h16e: qq = 8'h00; // 0x16e
	13'h16f: qq = 8'h00; // 0x16f
	13'h170: qq = 8'h00; // 0x170
	13'h171: qq = 8'h06; // 0x171
	13'h172: qq = 8'h06; // 0x172
	13'h173: qq = 8'h00; // 0x173
	13'h174: qq = 8'h00; // 0x174
	13'h175: qq = 8'h06; // 0x175
	13'h176: qq = 8'h06; // 0x176
	13'h177: qq = 8'h00; // 0x177
	13'h178: qq = 8'h00; // 0x178
	13'h179: qq = 8'h00; // 0x179
	13'h17a: qq = 8'h00; // 0x17a
	13'h17b: qq = 8'h00; // 0x17b
	13'h17c: qq = 8'h00; // 0x17c
	13'h17d: qq = 8'h06; // 0x17d
	13'h17e: qq = 8'h06; // 0x17e
	13'h17f: qq = 8'h00; // 0x17f
	13'h180: qq = 8'h00; // 0x180
	13'h181: qq = 8'h08; // 0x181
	13'h182: qq = 8'h0c; // 0x182
	13'h183: qq = 8'h06; // 0x183
	13'h184: qq = 8'h06; // 0x184
	13'h185: qq = 8'h06; // 0x185
	13'h186: qq = 8'h04; // 0x186
	13'h187: qq = 8'h08; // 0x187
	13'h188: qq = 8'h00; // 0x188
	13'h189: qq = 8'h00; // 0x189
	13'h18a: qq = 8'h00; // 0x18a
	13'h18b: qq = 8'h00; // 0x18b
	13'h18c: qq = 8'h00; // 0x18c
	13'h18d: qq = 8'h00; // 0x18d
	13'h18e: qq = 8'h00; // 0x18e
	13'h18f: qq = 8'h0c; // 0x18f
	13'h190: qq = 8'h00; // 0x190
	13'h191: qq = 8'h0c; // 0x191
	13'h192: qq = 8'h06; // 0x192
	13'h193: qq = 8'h0e; // 0x193
	13'h194: qq = 8'h0c; // 0x194
	13'h195: qq = 8'h08; // 0x195
	13'h196: qq = 8'h00; // 0x196
	13'h197: qq = 8'h0e; // 0x197
	13'h198: qq = 8'h00; // 0x198
	13'h199: qq = 8'h0e; // 0x199
	13'h19a: qq = 8'h0c; // 0x19a
	13'h19b: qq = 8'h08; // 0x19b
	13'h19c: qq = 8'h0c; // 0x19c
	13'h19d: qq = 8'h06; // 0x19d
	13'h19e: qq = 8'h06; // 0x19e
	13'h19f: qq = 8'h0c; // 0x19f
	13'h1a0: qq = 8'h00; // 0x1a0
	13'h1a1: qq = 8'h0c; // 0x1a1
	13'h1a2: qq = 8'h0c; // 0x1a2
	13'h1a3: qq = 8'h0c; // 0x1a3
	13'h1a4: qq = 8'h0c; // 0x1a4
	13'h1a5: qq = 8'h0e; // 0x1a5
	13'h1a6: qq = 8'h0c; // 0x1a6
	13'h1a7: qq = 8'h0c; // 0x1a7
	13'h1a8: qq = 8'h00; // 0x1a8
	13'h1a9: qq = 8'h0c; // 0x1a9
	13'h1aa: qq = 8'h00; // 0x1aa
	13'h1ab: qq = 8'h0c; // 0x1ab
	13'h1ac: qq = 8'h06; // 0x1ac
	13'h1ad: qq = 8'h06; // 0x1ad
	13'h1ae: qq = 8'h06; // 0x1ae
	13'h1af: qq = 8'h0c; // 0x1af
	13'h1b0: qq = 8'h00; // 0x1b0
	13'h1b1: qq = 8'h0c; // 0x1b1
	13'h1b2: qq = 8'h00; // 0x1b2
	13'h1b3: qq = 8'h00; // 0x1b3
	13'h1b4: qq = 8'h0c; // 0x1b4
	13'h1b5: qq = 8'h06; // 0x1b5
	13'h1b6: qq = 8'h06; // 0x1b6
	13'h1b7: qq = 8'h0c; // 0x1b7
	13'h1b8: qq = 8'h00; // 0x1b8
	13'h1b9: qq = 8'h0e; // 0x1b9
	13'h1ba: qq = 8'h06; // 0x1ba
	13'h1bb: qq = 8'h0c; // 0x1bb
	13'h1bc: qq = 8'h08; // 0x1bc
	13'h1bd: qq = 8'h00; // 0x1bd
	13'h1be: qq = 8'h00; // 0x1be
	13'h1bf: qq = 8'h00; // 0x1bf
	13'h1c0: qq = 8'h00; // 0x1c0
	13'h1c1: qq = 8'h08; // 0x1c1
	13'h1c2: qq = 8'h04; // 0x1c2
	13'h1c3: qq = 8'h04; // 0x1c3
	13'h1c4: qq = 8'h08; // 0x1c4
	13'h1c5: qq = 8'h0e; // 0x1c5
	13'h1c6: qq = 8'h06; // 0x1c6
	13'h1c7: qq = 8'h0c; // 0x1c7
	13'h1c8: qq = 8'h00; // 0x1c8
	13'h1c9: qq = 8'h0c; // 0x1c9
	13'h1ca: qq = 8'h06; // 0x1ca
	13'h1cb: qq = 8'h06; // 0x1cb
	13'h1cc: qq = 8'h0e; // 0x1cc
	13'h1cd: qq = 8'h06; // 0x1cd
	13'h1ce: qq = 8'h0c; // 0x1ce
	13'h1cf: qq = 8'h08; // 0x1cf
	13'h1d0: qq = 8'h00; // 0x1d0
	13'h1d1: qq = 8'h00; // 0x1d1
	13'h1d2: qq = 8'h00; // 0x1d2
	13'h1d3: qq = 8'h00; // 0x1d3
	13'h1d4: qq = 8'h00; // 0x1d4
	13'h1d5: qq = 8'h00; // 0x1d5
	13'h1d6: qq = 8'h00; // 0x1d6
	13'h1d7: qq = 8'h00; // 0x1d7
	13'h1d8: qq = 8'h00; // 0x1d8
	13'h1d9: qq = 8'h00; // 0x1d9
	13'h1da: qq = 8'h00; // 0x1da
	13'h1db: qq = 8'h00; // 0x1db
	13'h1dc: qq = 8'h00; // 0x1dc
	13'h1dd: qq = 8'h00; // 0x1dd
	13'h1de: qq = 8'h00; // 0x1de
	13'h1df: qq = 8'h00; // 0x1df
	13'h1e0: qq = 8'h00; // 0x1e0
	13'h1e1: qq = 8'h01; // 0x1e1
	13'h1e2: qq = 8'h07; // 0x1e2
	13'h1e3: qq = 8'h0f; // 0x1e3
	13'h1e4: qq = 8'h0f; // 0x1e4
	13'h1e5: qq = 8'h0f; // 0x1e5
	13'h1e6: qq = 8'h0f; // 0x1e6
	13'h1e7: qq = 8'h01; // 0x1e7
	13'h1e8: qq = 8'h00; // 0x1e8
	13'h1e9: qq = 8'h00; // 0x1e9
	13'h1ea: qq = 8'h00; // 0x1ea
	13'h1eb: qq = 8'h00; // 0x1eb
	13'h1ec: qq = 8'h0c; // 0x1ec
	13'h1ed: qq = 8'h0e; // 0x1ed
	13'h1ee: qq = 8'h0f; // 0x1ee
	13'h1ef: qq = 8'h0f; // 0x1ef
	13'h1f0: qq = 8'h05; // 0x1f0
	13'h1f1: qq = 8'h05; // 0x1f1
	13'h1f2: qq = 8'h01; // 0x1f2
	13'h1f3: qq = 8'h0f; // 0x1f3
	13'h1f4: qq = 8'h0f; // 0x1f4
	13'h1f5: qq = 8'h0f; // 0x1f5
	13'h1f6: qq = 8'h0f; // 0x1f6
	13'h1f7: qq = 8'h06; // 0x1f7
	13'h1f8: qq = 8'h0e; // 0x1f8
	13'h1f9: qq = 8'h06; // 0x1f9
	13'h1fa: qq = 8'h04; // 0x1fa
	13'h1fb: qq = 8'h0e; // 0x1fb
	13'h1fc: qq = 8'h0e; // 0x1fc
	13'h1fd: qq = 8'h0c; // 0x1fd
	13'h1fe: qq = 8'h08; // 0x1fe
	13'h1ff: qq = 8'h00; // 0x1ff
		endcase

	assign q = qq;
	endmodule // rom Char_MSB
